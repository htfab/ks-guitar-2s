magic
tech sky130A
magscale 1 2
timestamp 1641015008
<< locali >>
rect 102149 654211 102183 655265
rect 106657 654279 106691 655265
rect 115489 654551 115523 655265
rect 119905 654347 119939 655265
rect 128737 654415 128771 655265
rect 141801 654619 141835 655265
rect 146217 654823 146251 655265
rect 431141 654755 431175 654993
rect 448805 654687 448839 654993
rect 457453 654483 457487 654993
rect 488549 654143 488583 654993
rect 58541 50643 58575 50949
rect 63785 50847 63819 50949
rect 63693 50575 63727 50813
rect 67959 50677 68201 50711
rect 63785 50235 63819 50609
rect 81909 50099 81943 51017
rect 85589 51017 85865 51051
rect 85589 50983 85623 51017
rect 166089 50711 166123 50949
rect 173173 50847 173207 50949
rect 166215 50745 166365 50779
rect 88993 50507 89027 50677
rect 91143 50473 91293 50507
rect 97733 50371 97767 50473
rect 97825 50371 97859 50677
rect 173265 50643 173299 50949
rect 88993 50031 89027 50133
rect 125425 50031 125459 50337
rect 123895 49997 124079 50031
rect 89085 49827 89119 49997
rect 124045 49963 124079 49997
rect 153025 49895 153059 50541
rect 134383 49793 134625 49827
rect 172345 49759 172379 49929
rect 180533 49759 180567 50813
rect 533353 50507 533387 50813
rect 543013 50235 543047 50473
rect 50261 3451 50295 4029
rect 453865 3927 453899 4097
rect 548533 3927 548567 4029
rect 458373 3383 458407 3893
rect 548441 3451 548475 3893
rect 530501 2975 530535 3417
rect 552489 3179 552523 3417
rect 552581 3043 552615 3417
rect 552673 2907 552707 3009
<< viali >>
rect 102149 655265 102183 655299
rect 106657 655265 106691 655299
rect 115489 655265 115523 655299
rect 115489 654517 115523 654551
rect 119905 655265 119939 655299
rect 128737 655265 128771 655299
rect 141801 655265 141835 655299
rect 146217 655265 146251 655299
rect 146217 654789 146251 654823
rect 431141 654993 431175 655027
rect 431141 654721 431175 654755
rect 448805 654993 448839 655027
rect 448805 654653 448839 654687
rect 457453 654993 457487 655027
rect 141801 654585 141835 654619
rect 457453 654449 457487 654483
rect 488549 654993 488583 655027
rect 128737 654381 128771 654415
rect 119905 654313 119939 654347
rect 106657 654245 106691 654279
rect 102149 654177 102183 654211
rect 488549 654109 488583 654143
rect 81909 51017 81943 51051
rect 58541 50949 58575 50983
rect 63785 50949 63819 50983
rect 58541 50609 58575 50643
rect 63693 50813 63727 50847
rect 63785 50813 63819 50847
rect 67925 50677 67959 50711
rect 68201 50677 68235 50711
rect 63693 50541 63727 50575
rect 63785 50609 63819 50643
rect 63785 50201 63819 50235
rect 85865 51017 85899 51051
rect 85589 50949 85623 50983
rect 166089 50949 166123 50983
rect 173173 50949 173207 50983
rect 173173 50813 173207 50847
rect 173265 50949 173299 50983
rect 166181 50745 166215 50779
rect 166365 50745 166399 50779
rect 88993 50677 89027 50711
rect 97825 50677 97859 50711
rect 166089 50677 166123 50711
rect 88993 50473 89027 50507
rect 91109 50473 91143 50507
rect 91293 50473 91327 50507
rect 97733 50473 97767 50507
rect 97733 50337 97767 50371
rect 173265 50609 173299 50643
rect 180533 50813 180567 50847
rect 153025 50541 153059 50575
rect 97825 50337 97859 50371
rect 125425 50337 125459 50371
rect 81909 50065 81943 50099
rect 88993 50133 89027 50167
rect 88993 49997 89027 50031
rect 89085 49997 89119 50031
rect 123861 49997 123895 50031
rect 125425 49997 125459 50031
rect 124045 49929 124079 49963
rect 153025 49861 153059 49895
rect 172345 49929 172379 49963
rect 89085 49793 89119 49827
rect 134349 49793 134383 49827
rect 134625 49793 134659 49827
rect 172345 49725 172379 49759
rect 533353 50813 533387 50847
rect 533353 50473 533387 50507
rect 543013 50473 543047 50507
rect 543013 50201 543047 50235
rect 180533 49725 180567 49759
rect 453865 4097 453899 4131
rect 50261 4029 50295 4063
rect 548533 4029 548567 4063
rect 453865 3893 453899 3927
rect 458373 3893 458407 3927
rect 50261 3417 50295 3451
rect 548441 3893 548475 3927
rect 548533 3893 548567 3927
rect 458373 3349 458407 3383
rect 530501 3417 530535 3451
rect 548441 3417 548475 3451
rect 552489 3417 552523 3451
rect 552489 3145 552523 3179
rect 552581 3417 552615 3451
rect 552581 3009 552615 3043
rect 552673 3009 552707 3043
rect 530501 2941 530535 2975
rect 552673 2873 552707 2907
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 329834 700992 329840 701004
rect 154172 700964 329840 700992
rect 154172 700952 154178 700964
rect 329834 700952 329840 700964
rect 329892 700952 329898 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 325694 700924 325700 700936
rect 137888 700896 325700 700924
rect 137888 700884 137894 700896
rect 325694 700884 325700 700896
rect 325752 700884 325758 700936
rect 335998 700884 336004 700936
rect 336056 700924 336062 700936
rect 364978 700924 364984 700936
rect 336056 700896 364984 700924
rect 336056 700884 336062 700896
rect 364978 700884 364984 700896
rect 365036 700884 365042 700936
rect 260742 700816 260748 700868
rect 260800 700856 260806 700868
rect 462314 700856 462320 700868
rect 260800 700828 462320 700856
rect 260800 700816 260806 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 264882 700748 264888 700800
rect 264940 700788 264946 700800
rect 478506 700788 478512 700800
rect 264940 700760 478512 700788
rect 264940 700748 264946 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 343634 700720 343640 700732
rect 89220 700692 343640 700720
rect 89220 700680 89226 700692
rect 343634 700680 343640 700692
rect 343692 700680 343698 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 338114 700652 338120 700664
rect 73028 700624 338120 700652
rect 73028 700612 73034 700624
rect 338114 700612 338120 700624
rect 338172 700612 338178 700664
rect 340138 700612 340144 700664
rect 340196 700652 340202 700664
rect 494790 700652 494796 700664
rect 340196 700624 494796 700652
rect 340196 700612 340202 700624
rect 494790 700612 494796 700624
rect 494848 700612 494854 700664
rect 246942 700544 246948 700596
rect 247000 700584 247006 700596
rect 527174 700584 527180 700596
rect 247000 700556 527180 700584
rect 247000 700544 247006 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 252462 700476 252468 700528
rect 252520 700516 252526 700528
rect 543458 700516 543464 700528
rect 252520 700488 543464 700516
rect 252520 700476 252526 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 347774 700448 347780 700460
rect 40552 700420 347780 700448
rect 40552 700408 40558 700420
rect 347774 700408 347780 700420
rect 347832 700408 347838 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 356054 700380 356060 700392
rect 24360 700352 356060 700380
rect 24360 700340 24366 700352
rect 356054 700340 356060 700352
rect 356112 700340 356118 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 351914 700312 351920 700324
rect 8168 700284 351920 700312
rect 8168 700272 8174 700284
rect 351914 700272 351920 700284
rect 351972 700272 351978 700324
rect 542998 700272 543004 700324
rect 543056 700312 543062 700324
rect 559650 700312 559656 700324
rect 543056 700284 559656 700312
rect 543056 700272 543062 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 278682 700204 278688 700256
rect 278740 700244 278746 700256
rect 413646 700244 413652 700256
rect 278740 700216 413652 700244
rect 278740 700204 278746 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 274542 700136 274548 700188
rect 274600 700176 274606 700188
rect 397454 700176 397460 700188
rect 274600 700148 397460 700176
rect 274600 700136 274606 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 311894 700108 311900 700120
rect 202840 700080 311900 700108
rect 202840 700068 202846 700080
rect 311894 700068 311900 700080
rect 311952 700068 311958 700120
rect 218974 700000 218980 700052
rect 219032 700040 219038 700052
rect 316034 700040 316040 700052
rect 219032 700012 316040 700040
rect 219032 700000 219038 700012
rect 316034 700000 316040 700012
rect 316092 700000 316098 700052
rect 291102 699932 291108 699984
rect 291160 699972 291166 699984
rect 348786 699972 348792 699984
rect 291160 699944 348792 699972
rect 291160 699932 291166 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 286962 699864 286968 699916
rect 287020 699904 287026 699916
rect 332502 699904 332508 699916
rect 287020 699876 332508 699904
rect 287020 699864 287026 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 299566 699836 299572 699848
rect 267700 699808 299572 699836
rect 267700 699796 267706 699808
rect 299566 699796 299572 699808
rect 299624 699796 299630 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 303614 699768 303620 699780
rect 283892 699740 303620 699768
rect 283892 699728 283898 699740
rect 303614 699728 303620 699740
rect 303672 699728 303678 699780
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 173158 699700 173164 699712
rect 170364 699672 173164 699700
rect 170364 699660 170370 699672
rect 173158 699660 173164 699672
rect 173216 699660 173222 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 240778 699700 240784 699712
rect 235224 699672 240784 699700
rect 235224 699660 235230 699672
rect 240778 699660 240784 699672
rect 240836 699660 240842 699712
rect 296622 698912 296628 698964
rect 296680 698952 296686 698964
rect 300118 698952 300124 698964
rect 296680 698924 300124 698952
rect 296680 698912 296686 698924
rect 300118 698912 300124 698924
rect 300176 698912 300182 698964
rect 234522 696940 234528 696992
rect 234580 696980 234586 696992
rect 580166 696980 580172 696992
rect 234580 696952 580172 696980
rect 234580 696940 234586 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 238662 683204 238668 683256
rect 238720 683244 238726 683256
rect 580166 683244 580172 683256
rect 238720 683216 580172 683244
rect 238720 683204 238726 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 360194 683176 360200 683188
rect 3476 683148 360200 683176
rect 3476 683136 3482 683148
rect 360194 683136 360200 683148
rect 360252 683136 360258 683188
rect 229830 670760 229836 670812
rect 229888 670800 229894 670812
rect 580166 670800 580172 670812
rect 229888 670772 580172 670800
rect 229888 670760 229894 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 369854 670732 369860 670744
rect 3568 670704 369860 670732
rect 3568 670692 3574 670704
rect 369854 670692 369860 670704
rect 369912 670692 369918 670744
rect 282086 660288 282092 660340
rect 282144 660328 282150 660340
rect 335998 660328 336004 660340
rect 282144 660300 336004 660328
rect 282144 660288 282150 660300
rect 335998 660288 336004 660300
rect 336056 660288 336062 660340
rect 240778 659268 240784 659320
rect 240836 659308 240842 659320
rect 308490 659308 308496 659320
rect 240836 659280 308496 659308
rect 240836 659268 240842 659280
rect 308490 659268 308496 659280
rect 308548 659268 308554 659320
rect 255774 659200 255780 659252
rect 255832 659240 255838 659252
rect 340138 659240 340144 659252
rect 255832 659212 340144 659240
rect 255832 659200 255838 659212
rect 340138 659200 340144 659212
rect 340196 659200 340202 659252
rect 173158 659132 173164 659184
rect 173216 659172 173222 659184
rect 321646 659172 321652 659184
rect 173216 659144 321652 659172
rect 173216 659132 173222 659144
rect 321646 659132 321652 659144
rect 321704 659132 321710 659184
rect 268930 659064 268936 659116
rect 268988 659104 268994 659116
rect 429194 659104 429200 659116
rect 268988 659076 429200 659104
rect 268988 659064 268994 659076
rect 429194 659064 429200 659076
rect 429252 659064 429258 659116
rect 106182 658996 106188 659048
rect 106240 659036 106246 659048
rect 334802 659036 334808 659048
rect 106240 659008 334808 659036
rect 106240 658996 106246 659008
rect 334802 658996 334808 659008
rect 334860 658996 334866 659048
rect 242526 658928 242532 658980
rect 242584 658968 242590 658980
rect 542998 658968 543004 658980
rect 242584 658940 543004 658968
rect 242584 658928 242590 658940
rect 542998 658928 543004 658940
rect 543056 658928 543062 658980
rect 29638 658316 29644 658368
rect 29696 658356 29702 658368
rect 541342 658356 541348 658368
rect 29696 658328 541348 658356
rect 29696 658316 29702 658328
rect 541342 658316 541348 658328
rect 541400 658316 541406 658368
rect 53650 658248 53656 658300
rect 53708 658288 53714 658300
rect 566458 658288 566464 658300
rect 53708 658260 566464 658288
rect 53708 658248 53714 658260
rect 566458 658248 566464 658260
rect 566516 658248 566522 658300
rect 211798 658180 211804 658232
rect 211856 658220 211862 658232
rect 565170 658220 565176 658232
rect 211856 658192 565176 658220
rect 211856 658180 211862 658192
rect 565170 658180 565176 658192
rect 565228 658180 565234 658232
rect 194226 658112 194232 658164
rect 194284 658152 194290 658164
rect 548610 658152 548616 658164
rect 194284 658124 548616 658152
rect 194284 658112 194290 658124
rect 548610 658112 548616 658124
rect 548668 658112 548674 658164
rect 3418 658044 3424 658096
rect 3476 658084 3482 658096
rect 365622 658084 365628 658096
rect 3476 658056 365628 658084
rect 3476 658044 3482 658056
rect 365622 658044 365628 658056
rect 365680 658044 365686 658096
rect 42242 657976 42248 658028
rect 42300 658016 42306 658028
rect 409506 658016 409512 658028
rect 42300 657988 409512 658016
rect 42300 657976 42306 657988
rect 409506 657976 409512 657988
rect 409564 657976 409570 658028
rect 132770 657908 132776 657960
rect 132828 657948 132834 657960
rect 184842 657948 184848 657960
rect 132828 657920 184848 657948
rect 132828 657908 132834 657920
rect 184842 657908 184848 657920
rect 184900 657908 184906 657960
rect 185486 657908 185492 657960
rect 185544 657948 185550 657960
rect 556890 657948 556896 657960
rect 185544 657920 556896 657948
rect 185544 657908 185550 657920
rect 556890 657908 556896 657920
rect 556948 657908 556954 657960
rect 167914 657840 167920 657892
rect 167972 657880 167978 657892
rect 551370 657880 551376 657892
rect 167972 657852 551376 657880
rect 167972 657840 167978 657852
rect 551370 657840 551376 657852
rect 551428 657840 551434 657892
rect 181070 657772 181076 657824
rect 181128 657812 181134 657824
rect 576210 657812 576216 657824
rect 181128 657784 576216 657812
rect 181128 657772 181134 657784
rect 576210 657772 576216 657784
rect 576268 657772 576274 657824
rect 25590 657704 25596 657756
rect 25648 657744 25654 657756
rect 435910 657744 435916 657756
rect 25648 657716 435916 657744
rect 25648 657704 25654 657716
rect 435910 657704 435916 657716
rect 435968 657704 435974 657756
rect 163498 657636 163504 657688
rect 163556 657676 163562 657688
rect 573450 657676 573456 657688
rect 163556 657648 573456 657676
rect 163556 657636 163562 657648
rect 573450 657636 573456 657648
rect 573508 657636 573514 657688
rect 154666 657568 154672 657620
rect 154724 657608 154730 657620
rect 574830 657608 574836 657620
rect 154724 657580 574836 657608
rect 154724 657568 154730 657580
rect 574830 657568 574836 657580
rect 574888 657568 574894 657620
rect 137094 657500 137100 657552
rect 137152 657540 137158 657552
rect 566550 657540 566556 657552
rect 137152 657512 566556 657540
rect 137152 657500 137158 657512
rect 566550 657500 566556 657512
rect 566608 657500 566614 657552
rect 39298 657432 39304 657484
rect 39356 657472 39362 657484
rect 471054 657472 471060 657484
rect 39356 657444 471060 657472
rect 39356 657432 39362 657444
rect 471054 657432 471060 657444
rect 471112 657432 471118 657484
rect 36538 657364 36544 657416
rect 36596 657404 36602 657416
rect 475378 657404 475384 657416
rect 36596 657376 475384 657404
rect 36596 657364 36602 657376
rect 475378 657364 475384 657376
rect 475436 657364 475442 657416
rect 11698 657296 11704 657348
rect 11756 657336 11762 657348
rect 462222 657336 462228 657348
rect 11756 657308 462228 657336
rect 11756 657296 11762 657308
rect 462222 657296 462228 657308
rect 462280 657296 462286 657348
rect 110782 657228 110788 657280
rect 110840 657268 110846 657280
rect 562410 657268 562416 657280
rect 110840 657240 562416 657268
rect 110840 657228 110846 657240
rect 562410 657228 562416 657240
rect 562468 657228 562474 657280
rect 42058 657160 42064 657212
rect 42116 657200 42122 657212
rect 501782 657200 501788 657212
rect 42116 657172 501788 657200
rect 42116 657160 42122 657172
rect 501782 657160 501788 657172
rect 501840 657160 501846 657212
rect 88794 657092 88800 657144
rect 88852 657132 88858 657144
rect 548518 657132 548524 657144
rect 88852 657104 548524 657132
rect 88852 657092 88858 657104
rect 548518 657092 548524 657104
rect 548576 657092 548582 657144
rect 15838 657024 15844 657076
rect 15896 657064 15902 657076
rect 484210 657064 484216 657076
rect 15896 657036 484216 657064
rect 15896 657024 15902 657036
rect 484210 657024 484216 657036
rect 484268 657024 484274 657076
rect 75638 656956 75644 657008
rect 75696 656996 75702 657008
rect 545758 656996 545764 657008
rect 75696 656968 545764 656996
rect 75696 656956 75702 656968
rect 545758 656956 545764 656968
rect 545816 656956 545822 657008
rect 84378 656888 84384 656940
rect 84436 656928 84442 656940
rect 558178 656928 558184 656940
rect 84436 656900 558184 656928
rect 84436 656888 84442 656900
rect 558178 656888 558184 656900
rect 558236 656888 558242 656940
rect 216214 656820 216220 656872
rect 216272 656860 216278 656872
rect 548702 656860 548708 656872
rect 216272 656832 548708 656860
rect 216272 656820 216278 656832
rect 548702 656820 548708 656832
rect 548760 656820 548766 656872
rect 203058 656752 203064 656804
rect 203116 656792 203122 656804
rect 547230 656792 547236 656804
rect 203116 656764 547236 656792
rect 203116 656752 203122 656764
rect 547230 656752 547236 656764
rect 547288 656752 547294 656804
rect 189810 656684 189816 656736
rect 189868 656724 189874 656736
rect 545850 656724 545856 656736
rect 189868 656696 545856 656724
rect 189868 656684 189874 656696
rect 545850 656684 545856 656696
rect 545908 656684 545914 656736
rect 11882 656616 11888 656668
rect 11940 656656 11946 656668
rect 374362 656656 374368 656668
rect 11940 656628 374368 656656
rect 11940 656616 11946 656628
rect 374362 656616 374368 656628
rect 374420 656616 374426 656668
rect 176654 656548 176660 656600
rect 176712 656588 176718 656600
rect 544470 656588 544476 656600
rect 176712 656560 544476 656588
rect 176712 656548 176718 656560
rect 544470 656548 544476 656560
rect 544528 656548 544534 656600
rect 14550 656480 14556 656532
rect 14608 656520 14614 656532
rect 387518 656520 387524 656532
rect 14608 656492 387524 656520
rect 14608 656480 14614 656492
rect 387518 656480 387524 656492
rect 387576 656480 387582 656532
rect 15930 656412 15936 656464
rect 15988 656452 15994 656464
rect 400766 656452 400772 656464
rect 15988 656424 400772 656452
rect 15988 656412 15994 656424
rect 400766 656412 400772 656424
rect 400824 656412 400830 656464
rect 17310 656344 17316 656396
rect 17368 656384 17374 656396
rect 413922 656384 413928 656396
rect 17368 656356 413928 656384
rect 17368 656344 17374 656356
rect 413922 656344 413928 656356
rect 413980 656344 413986 656396
rect 159082 656276 159088 656328
rect 159140 656316 159146 656328
rect 555510 656316 555516 656328
rect 159140 656288 555516 656316
rect 159140 656276 159146 656288
rect 555510 656276 555516 656288
rect 555568 656276 555574 656328
rect 18690 656208 18696 656260
rect 18748 656248 18754 656260
rect 427078 656248 427084 656260
rect 18748 656220 427084 656248
rect 18748 656208 18754 656220
rect 427078 656208 427084 656220
rect 427136 656208 427142 656260
rect 172238 656140 172244 656192
rect 172296 656180 172302 656192
rect 580350 656180 580356 656192
rect 172296 656152 580356 656180
rect 172296 656140 172302 656152
rect 580350 656140 580356 656152
rect 580408 656140 580414 656192
rect 21450 656072 21456 656124
rect 21508 656112 21514 656124
rect 440234 656112 440240 656124
rect 21508 656084 440240 656112
rect 21508 656072 21514 656084
rect 440234 656072 440240 656084
rect 440292 656072 440298 656124
rect 22738 656004 22744 656056
rect 22796 656044 22802 656056
rect 453482 656044 453488 656056
rect 22796 656016 453488 656044
rect 22796 656004 22802 656016
rect 453482 656004 453488 656016
rect 453540 656004 453546 656056
rect 25498 655936 25504 655988
rect 25556 655976 25562 655988
rect 466638 655976 466644 655988
rect 25556 655948 466644 655976
rect 25556 655936 25562 655948
rect 466638 655936 466644 655948
rect 466696 655936 466702 655988
rect 123938 655868 123944 655920
rect 123996 655908 124002 655920
rect 565078 655908 565084 655920
rect 123996 655880 565084 655908
rect 123996 655868 124002 655880
rect 565078 655868 565084 655880
rect 565136 655868 565142 655920
rect 29730 655800 29736 655852
rect 29788 655840 29794 655852
rect 492950 655840 492956 655852
rect 29788 655812 492956 655840
rect 29788 655800 29794 655812
rect 492950 655800 492956 655812
rect 493008 655800 493014 655852
rect 97626 655732 97632 655784
rect 97684 655772 97690 655784
rect 561030 655772 561036 655784
rect 97684 655744 561036 655772
rect 97684 655732 97690 655744
rect 561030 655732 561036 655744
rect 561088 655732 561094 655784
rect 7558 655664 7564 655716
rect 7616 655704 7622 655716
rect 479518 655704 479524 655716
rect 7616 655676 479524 655704
rect 7616 655664 7622 655676
rect 479518 655664 479524 655676
rect 479576 655664 479582 655716
rect 32398 655596 32404 655648
rect 32456 655636 32462 655648
rect 505830 655636 505836 655648
rect 32456 655608 505836 655636
rect 32456 655596 32462 655608
rect 505830 655596 505836 655608
rect 505888 655596 505894 655648
rect 71498 655528 71504 655580
rect 71556 655568 71562 655580
rect 556798 655568 556804 655580
rect 71556 655540 556804 655568
rect 71556 655528 71562 655540
rect 556798 655528 556804 655540
rect 556856 655528 556862 655580
rect 184842 655392 184848 655444
rect 184900 655432 184906 655444
rect 580258 655432 580264 655444
rect 184900 655404 580264 655432
rect 184900 655392 184906 655404
rect 580258 655392 580264 655404
rect 580316 655392 580322 655444
rect 225322 655324 225328 655376
rect 225380 655364 225386 655376
rect 558362 655364 558368 655376
rect 225380 655336 558368 655364
rect 225380 655324 225386 655336
rect 558362 655324 558368 655336
rect 558420 655324 558426 655376
rect 102134 655296 102140 655308
rect 102095 655268 102140 655296
rect 102134 655256 102140 655268
rect 102192 655256 102198 655308
rect 106642 655296 106648 655308
rect 106603 655268 106648 655296
rect 106642 655256 106648 655268
rect 106700 655256 106706 655308
rect 115474 655296 115480 655308
rect 115435 655268 115480 655296
rect 115474 655256 115480 655268
rect 115532 655256 115538 655308
rect 119890 655296 119896 655308
rect 119851 655268 119896 655296
rect 119890 655256 119896 655268
rect 119948 655256 119954 655308
rect 128722 655296 128728 655308
rect 128683 655268 128728 655296
rect 128722 655256 128728 655268
rect 128780 655256 128786 655308
rect 141786 655296 141792 655308
rect 141747 655268 141792 655296
rect 141786 655256 141792 655268
rect 141844 655256 141850 655308
rect 146202 655296 146208 655308
rect 146163 655268 146208 655296
rect 146202 655256 146208 655268
rect 146260 655256 146266 655308
rect 198550 655256 198556 655308
rect 198608 655296 198614 655308
rect 554038 655296 554044 655308
rect 198608 655268 554044 655296
rect 198608 655256 198614 655268
rect 554038 655256 554044 655268
rect 554096 655256 554102 655308
rect 40770 655188 40776 655240
rect 40828 655228 40834 655240
rect 404814 655228 404820 655240
rect 40828 655200 404820 655228
rect 40828 655188 40834 655200
rect 404814 655188 404820 655200
rect 404872 655188 404878 655240
rect 7650 655120 7656 655172
rect 7708 655160 7714 655172
rect 382918 655160 382924 655172
rect 7708 655132 382924 655160
rect 7708 655120 7714 655132
rect 382918 655120 382924 655132
rect 382976 655120 382982 655172
rect 42150 655052 42156 655104
rect 42208 655092 42214 655104
rect 418154 655092 418160 655104
rect 42208 655064 418160 655092
rect 42208 655052 42214 655064
rect 418154 655052 418160 655064
rect 418212 655052 418218 655104
rect 10318 654984 10324 655036
rect 10376 655024 10382 655036
rect 396074 655024 396080 655036
rect 10376 654996 396080 655024
rect 10376 654984 10382 654996
rect 396074 654984 396080 654996
rect 396132 654984 396138 655036
rect 422478 655024 422484 655036
rect 412606 654996 422484 655024
rect 22830 654916 22836 654968
rect 22888 654956 22894 654968
rect 412606 654956 412634 654996
rect 422478 654984 422484 654996
rect 422536 654984 422542 655036
rect 431126 655024 431132 655036
rect 431087 654996 431132 655024
rect 431126 654984 431132 654996
rect 431184 654984 431190 655036
rect 444374 654984 444380 655036
rect 444432 654984 444438 655036
rect 448790 655024 448796 655036
rect 448751 654996 448796 655024
rect 448790 654984 448796 654996
rect 448848 654984 448854 655036
rect 457438 655024 457444 655036
rect 457399 654996 457444 655024
rect 457438 654984 457444 654996
rect 457496 654984 457502 655036
rect 488534 655024 488540 655036
rect 488495 654996 488540 655024
rect 488534 654984 488540 654996
rect 488592 654984 488598 655036
rect 22888 654928 412634 654956
rect 22888 654916 22894 654928
rect 36630 654848 36636 654900
rect 36688 654888 36694 654900
rect 444392 654888 444420 654984
rect 36688 654860 444420 654888
rect 36688 654848 36694 654860
rect 146205 654823 146263 654829
rect 146205 654789 146217 654823
rect 146251 654820 146263 654823
rect 558270 654820 558276 654832
rect 146251 654792 558276 654820
rect 146251 654789 146263 654792
rect 146205 654783 146263 654789
rect 558270 654780 558276 654792
rect 558328 654780 558334 654832
rect 11790 654712 11796 654764
rect 11848 654752 11854 654764
rect 431129 654755 431187 654761
rect 431129 654752 431141 654755
rect 11848 654724 431141 654752
rect 11848 654712 11854 654724
rect 431129 654721 431141 654724
rect 431175 654721 431187 654755
rect 431129 654715 431187 654721
rect 26878 654644 26884 654696
rect 26936 654684 26942 654696
rect 448793 654687 448851 654693
rect 448793 654684 448805 654687
rect 26936 654656 448805 654684
rect 26936 654644 26942 654656
rect 448793 654653 448805 654656
rect 448839 654653 448851 654687
rect 448793 654647 448851 654653
rect 141789 654619 141847 654625
rect 141789 654585 141801 654619
rect 141835 654616 141847 654619
rect 569218 654616 569224 654628
rect 141835 654588 569224 654616
rect 141835 654585 141847 654588
rect 141789 654579 141847 654585
rect 569218 654576 569224 654588
rect 569276 654576 569282 654628
rect 115477 654551 115535 654557
rect 115477 654517 115489 654551
rect 115523 654548 115535 654551
rect 544378 654548 544384 654560
rect 115523 654520 544384 654548
rect 115523 654517 115535 654520
rect 115477 654511 115535 654517
rect 544378 654508 544384 654520
rect 544436 654508 544442 654560
rect 14458 654440 14464 654492
rect 14516 654480 14522 654492
rect 457441 654483 457499 654489
rect 457441 654480 457453 654483
rect 14516 654452 457453 654480
rect 14516 654440 14522 654452
rect 457441 654449 457453 654452
rect 457487 654449 457499 654483
rect 457441 654443 457499 654449
rect 128725 654415 128783 654421
rect 128725 654381 128737 654415
rect 128771 654412 128783 654415
rect 573358 654412 573364 654424
rect 128771 654384 573364 654412
rect 128771 654381 128783 654384
rect 128725 654375 128783 654381
rect 573358 654372 573364 654384
rect 573416 654372 573422 654424
rect 119893 654347 119951 654353
rect 119893 654313 119905 654347
rect 119939 654344 119951 654347
rect 578878 654344 578884 654356
rect 119939 654316 578884 654344
rect 119939 654313 119951 654316
rect 119893 654307 119951 654313
rect 578878 654304 578884 654316
rect 578936 654304 578942 654356
rect 106645 654279 106703 654285
rect 106645 654245 106657 654279
rect 106691 654276 106703 654279
rect 571978 654276 571984 654288
rect 106691 654248 571984 654276
rect 106691 654245 106703 654248
rect 106645 654239 106703 654245
rect 571978 654236 571984 654248
rect 572036 654236 572042 654288
rect 102137 654211 102195 654217
rect 102137 654177 102149 654211
rect 102183 654208 102195 654211
rect 576118 654208 576124 654220
rect 102183 654180 576124 654208
rect 102183 654177 102195 654180
rect 102137 654171 102195 654177
rect 576118 654168 576124 654180
rect 576176 654168 576182 654220
rect 3510 654100 3516 654152
rect 3568 654140 3574 654152
rect 488537 654143 488595 654149
rect 488537 654140 488549 654143
rect 3568 654112 488549 654140
rect 3568 654100 3574 654112
rect 488537 654109 488549 654112
rect 488583 654109 488595 654143
rect 488537 654103 488595 654109
rect 561122 644376 561128 644428
rect 561180 644416 561186 644428
rect 580166 644416 580172 644428
rect 561180 644388 580172 644416
rect 561180 644376 561186 644388
rect 580166 644376 580172 644388
rect 580224 644376 580230 644428
rect 3326 633360 3332 633412
rect 3384 633400 3390 633412
rect 11882 633400 11888 633412
rect 3384 633372 11888 633400
rect 3384 633360 3390 633372
rect 11882 633360 11888 633372
rect 11940 633360 11946 633412
rect 558362 632000 558368 632052
rect 558420 632040 558426 632052
rect 580166 632040 580172 632052
rect 558420 632012 580172 632040
rect 558420 632000 558426 632012
rect 580166 632000 580172 632012
rect 580224 632000 580230 632052
rect 3142 619284 3148 619336
rect 3200 619324 3206 619336
rect 7650 619324 7656 619336
rect 3200 619296 7656 619324
rect 3200 619284 3206 619296
rect 7650 619284 7656 619296
rect 7708 619284 7714 619336
rect 548702 618196 548708 618248
rect 548760 618236 548766 618248
rect 580166 618236 580172 618248
rect 548760 618208 580172 618236
rect 548760 618196 548766 618208
rect 580166 618196 580172 618208
rect 580224 618196 580230 618248
rect 3050 607112 3056 607164
rect 3108 607152 3114 607164
rect 36722 607152 36728 607164
rect 3108 607124 36728 607152
rect 3108 607112 3114 607124
rect 36722 607112 36728 607124
rect 36780 607112 36786 607164
rect 555602 591948 555608 592000
rect 555660 591988 555666 592000
rect 580166 591988 580172 592000
rect 555660 591960 580172 591988
rect 555660 591948 555666 591960
rect 580166 591948 580172 591960
rect 580224 591948 580230 592000
rect 3326 580932 3332 580984
rect 3384 580972 3390 580984
rect 14550 580972 14556 580984
rect 3384 580944 14556 580972
rect 3384 580932 3390 580944
rect 14550 580932 14556 580944
rect 14608 580932 14614 580984
rect 565170 578144 565176 578196
rect 565228 578184 565234 578196
rect 579614 578184 579620 578196
rect 565228 578156 579620 578184
rect 565228 578144 565234 578156
rect 579614 578144 579620 578156
rect 579672 578144 579678 578196
rect 3326 567128 3332 567180
rect 3384 567168 3390 567180
rect 10318 567168 10324 567180
rect 3384 567140 10324 567168
rect 3384 567128 3390 567140
rect 10318 567128 10324 567140
rect 10376 567128 10382 567180
rect 547230 564340 547236 564392
rect 547288 564380 547294 564392
rect 580166 564380 580172 564392
rect 547288 564352 580172 564380
rect 547288 564340 547294 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 3326 554684 3332 554736
rect 3384 554724 3390 554736
rect 39390 554724 39396 554736
rect 3384 554696 39396 554724
rect 3384 554684 3390 554696
rect 39390 554684 39396 554696
rect 39448 554684 39454 554736
rect 548610 538160 548616 538212
rect 548668 538200 548674 538212
rect 580166 538200 580172 538212
rect 548668 538172 580172 538200
rect 548668 538160 548674 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 3326 528504 3332 528556
rect 3384 528544 3390 528556
rect 15930 528544 15936 528556
rect 3384 528516 15936 528544
rect 3384 528504 3390 528516
rect 15930 528504 15936 528516
rect 15988 528504 15994 528556
rect 554038 525716 554044 525768
rect 554096 525756 554102 525768
rect 579890 525756 579896 525768
rect 554096 525728 579896 525756
rect 554096 525716 554102 525728
rect 579890 525716 579896 525728
rect 579948 525716 579954 525768
rect 3142 516060 3148 516112
rect 3200 516100 3206 516112
rect 42242 516100 42248 516112
rect 3200 516072 42248 516100
rect 3200 516060 3206 516072
rect 42242 516060 42248 516072
rect 42300 516060 42306 516112
rect 545850 511912 545856 511964
rect 545908 511952 545914 511964
rect 580166 511952 580172 511964
rect 545908 511924 580172 511952
rect 545908 511912 545914 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 2958 502256 2964 502308
rect 3016 502296 3022 502308
rect 40770 502296 40776 502308
rect 3016 502268 40776 502296
rect 3016 502256 3022 502268
rect 40770 502256 40776 502268
rect 40828 502256 40834 502308
rect 576210 485732 576216 485784
rect 576268 485772 576274 485784
rect 580166 485772 580172 485784
rect 576268 485744 580172 485772
rect 576268 485732 576274 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 3234 476008 3240 476060
rect 3292 476048 3298 476060
rect 17310 476048 17316 476060
rect 3292 476020 17316 476048
rect 3292 476008 3298 476020
rect 17310 476008 17316 476020
rect 17368 476008 17374 476060
rect 556890 471928 556896 471980
rect 556948 471968 556954 471980
rect 579614 471968 579620 471980
rect 556948 471940 579620 471968
rect 556948 471928 556954 471940
rect 579614 471928 579620 471940
rect 579672 471928 579678 471980
rect 3050 463632 3056 463684
rect 3108 463672 3114 463684
rect 22830 463672 22836 463684
rect 3108 463644 22836 463672
rect 3108 463632 3114 463644
rect 22830 463632 22836 463644
rect 22888 463632 22894 463684
rect 544470 458124 544476 458176
rect 544528 458164 544534 458176
rect 580166 458164 580172 458176
rect 544528 458136 580172 458164
rect 544528 458124 544534 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 42150 449868 42156 449880
rect 3384 449840 42156 449868
rect 3384 449828 3390 449840
rect 42150 449828 42156 449840
rect 42208 449828 42214 449880
rect 551370 431876 551376 431928
rect 551428 431916 551434 431928
rect 579614 431916 579620 431928
rect 551428 431888 579620 431916
rect 551428 431876 551434 431888
rect 579614 431876 579620 431888
rect 579672 431876 579678 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 18690 423620 18696 423632
rect 3384 423592 18696 423620
rect 3384 423580 3390 423592
rect 18690 423580 18696 423592
rect 18748 423580 18754 423632
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 25590 411244 25596 411256
rect 3016 411216 25596 411244
rect 3016 411204 3022 411216
rect 25590 411204 25596 411216
rect 25648 411204 25654 411256
rect 573450 405628 573456 405680
rect 573508 405668 573514 405680
rect 579614 405668 579620 405680
rect 573508 405640 579620 405668
rect 573508 405628 573514 405640
rect 579614 405628 579620 405640
rect 579672 405628 579678 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 11790 398800 11796 398812
rect 3384 398772 11796 398800
rect 3384 398760 3390 398772
rect 11790 398760 11796 398772
rect 11848 398760 11854 398812
rect 574830 379448 574836 379500
rect 574888 379488 574894 379500
rect 580166 379488 580172 379500
rect 574888 379460 580172 379488
rect 574888 379448 574894 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 21450 372552 21456 372564
rect 3384 372524 21456 372552
rect 3384 372512 3390 372524
rect 21450 372512 21456 372524
rect 21508 372512 21514 372564
rect 555510 365644 555516 365696
rect 555568 365684 555574 365696
rect 580166 365684 580172 365696
rect 555568 365656 580172 365684
rect 555568 365644 555574 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 26878 358748 26884 358760
rect 3384 358720 26884 358748
rect 3384 358708 3390 358720
rect 26878 358708 26884 358720
rect 26936 358708 26942 358760
rect 569310 353200 569316 353252
rect 569368 353240 569374 353252
rect 580166 353240 580172 353252
rect 569368 353212 580172 353240
rect 569368 353200 569374 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 36630 346372 36636 346384
rect 3384 346344 36636 346372
rect 3384 346332 3390 346344
rect 36630 346332 36636 346344
rect 36688 346332 36694 346384
rect 569218 325592 569224 325644
rect 569276 325632 569282 325644
rect 579890 325632 579896 325644
rect 569276 325604 579896 325632
rect 569276 325592 569282 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 22738 320124 22744 320136
rect 3384 320096 22744 320124
rect 3384 320084 3390 320096
rect 22738 320084 22744 320096
rect 22796 320084 22802 320136
rect 558270 313216 558276 313268
rect 558328 313256 558334 313268
rect 580166 313256 580172 313268
rect 558328 313228 580172 313256
rect 558328 313216 558334 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 11698 306320 11704 306332
rect 3384 306292 11704 306320
rect 3384 306280 3390 306292
rect 11698 306280 11704 306292
rect 11756 306280 11762 306332
rect 566550 299412 566556 299464
rect 566608 299452 566614 299464
rect 579614 299452 579620 299464
rect 566608 299424 579620 299452
rect 566608 299412 566614 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 3326 293904 3332 293956
rect 3384 293944 3390 293956
rect 14458 293944 14464 293956
rect 3384 293916 14464 293944
rect 3384 293904 3390 293916
rect 14458 293904 14464 293916
rect 14516 293904 14522 293956
rect 573358 273164 573364 273216
rect 573416 273204 573422 273216
rect 579890 273204 579896 273216
rect 573416 273176 579896 273204
rect 573416 273164 573422 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 25498 267696 25504 267708
rect 3016 267668 25504 267696
rect 3016 267656 3022 267668
rect 25498 267656 25504 267668
rect 25556 267656 25562 267708
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 36538 255252 36544 255264
rect 3200 255224 36544 255252
rect 3200 255212 3206 255224
rect 36538 255212 36544 255224
rect 36596 255212 36602 255264
rect 565078 245556 565084 245608
rect 565136 245596 565142 245608
rect 580166 245596 580172 245608
rect 565136 245568 580172 245596
rect 565136 245556 565142 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 39298 241448 39304 241460
rect 3292 241420 39304 241448
rect 3292 241408 3298 241420
rect 39298 241408 39304 241420
rect 39356 241408 39362 241460
rect 544378 233180 544384 233232
rect 544436 233220 544442 233232
rect 579982 233220 579988 233232
rect 544436 233192 579988 233220
rect 544436 233180 544442 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 3326 214956 3332 215008
rect 3384 214996 3390 215008
rect 7558 214996 7564 215008
rect 3384 214968 7564 214996
rect 3384 214956 3390 214968
rect 7558 214956 7564 214968
rect 7616 214956 7622 215008
rect 562410 206932 562416 206984
rect 562468 206972 562474 206984
rect 579798 206972 579804 206984
rect 562468 206944 579804 206972
rect 562468 206932 562474 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 576118 193128 576124 193180
rect 576176 193168 576182 193180
rect 580166 193168 580172 193180
rect 576176 193140 580172 193168
rect 576176 193128 576182 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 15838 189020 15844 189032
rect 3568 188992 15844 189020
rect 3568 188980 3574 188992
rect 15838 188980 15844 188992
rect 15896 188980 15902 189032
rect 571978 179324 571984 179376
rect 572036 179364 572042 179376
rect 580166 179364 580172 179376
rect 572036 179336 580172 179364
rect 572036 179324 572042 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 561030 166948 561036 167000
rect 561088 166988 561094 167000
rect 580166 166988 580172 167000
rect 561088 166960 580172 166988
rect 561088 166948 561094 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 29730 164200 29736 164212
rect 3292 164172 29736 164200
rect 3292 164160 3298 164172
rect 29730 164160 29736 164172
rect 29788 164160 29794 164212
rect 548518 153144 548524 153196
rect 548576 153184 548582 153196
rect 580166 153184 580172 153196
rect 548576 153156 580172 153184
rect 548576 153144 548582 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 42058 150396 42064 150408
rect 3568 150368 42064 150396
rect 3568 150356 3574 150368
rect 42058 150356 42064 150368
rect 42116 150356 42122 150408
rect 570598 139340 570604 139392
rect 570656 139380 570662 139392
rect 580166 139380 580172 139392
rect 570656 139352 580172 139380
rect 570656 139340 570662 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 40678 137952 40684 137964
rect 3568 137924 40684 137952
rect 3568 137912 3574 137924
rect 40678 137912 40684 137924
rect 40736 137912 40742 137964
rect 558178 126896 558184 126948
rect 558236 126936 558242 126948
rect 580166 126936 580172 126948
rect 558236 126908 580172 126936
rect 558236 126896 558242 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 545758 113092 545764 113144
rect 545816 113132 545822 113144
rect 579798 113132 579804 113144
rect 545816 113104 579804 113132
rect 545816 113092 545822 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 32398 111772 32404 111784
rect 3200 111744 32404 111772
rect 3200 111732 3206 111744
rect 32398 111732 32404 111744
rect 32456 111732 32462 111784
rect 560938 100648 560944 100700
rect 560996 100688 561002 100700
rect 580166 100688 580172 100700
rect 560996 100660 580172 100688
rect 560996 100648 561002 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 556798 86912 556804 86964
rect 556856 86952 556862 86964
rect 580166 86952 580172 86964
rect 556856 86924 580172 86952
rect 556856 86912 556862 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 17218 85524 17224 85536
rect 3200 85496 17224 85524
rect 3200 85484 3206 85496
rect 17218 85484 17224 85496
rect 17276 85484 17282 85536
rect 547138 73108 547144 73160
rect 547196 73148 547202 73160
rect 580166 73148 580172 73160
rect 547196 73120 580172 73148
rect 547196 73108 547202 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 33778 71720 33784 71732
rect 3476 71692 33784 71720
rect 3476 71680 3482 71692
rect 33778 71680 33784 71692
rect 33836 71680 33842 71732
rect 562318 60664 562324 60716
rect 562376 60704 562382 60716
rect 580166 60704 580172 60716
rect 562376 60676 580172 60704
rect 562376 60664 562382 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 2774 58624 2780 58676
rect 2832 58664 2838 58676
rect 4798 58664 4804 58676
rect 2832 58636 4804 58664
rect 2832 58624 2838 58636
rect 4798 58624 4804 58636
rect 4856 58624 4862 58676
rect 85408 51088 85804 51116
rect 23382 51008 23388 51060
rect 23440 51048 23446 51060
rect 62482 51048 62488 51060
rect 23440 51020 62488 51048
rect 23440 51008 23446 51020
rect 62482 51008 62488 51020
rect 62540 51008 62546 51060
rect 71038 51008 71044 51060
rect 71096 51048 71102 51060
rect 81802 51048 81808 51060
rect 71096 51020 81808 51048
rect 71096 51008 71102 51020
rect 81802 51008 81808 51020
rect 81860 51008 81866 51060
rect 81897 51051 81955 51057
rect 81897 51017 81909 51051
rect 81943 51048 81955 51051
rect 85408 51048 85436 51088
rect 81943 51020 85436 51048
rect 81943 51017 81955 51020
rect 81897 51011 81955 51017
rect 19242 50940 19248 50992
rect 19300 50980 19306 50992
rect 58434 50980 58440 50992
rect 19300 50952 58440 50980
rect 19300 50940 19306 50952
rect 58434 50940 58440 50952
rect 58492 50940 58498 50992
rect 58529 50983 58587 50989
rect 58529 50949 58541 50983
rect 58575 50980 58587 50983
rect 63773 50983 63831 50989
rect 63773 50980 63785 50983
rect 58575 50952 63785 50980
rect 58575 50949 58587 50952
rect 58529 50943 58587 50949
rect 63773 50949 63785 50952
rect 63819 50949 63831 50983
rect 78766 50980 78772 50992
rect 63773 50943 63831 50949
rect 64846 50952 78772 50980
rect 16482 50872 16488 50924
rect 16540 50912 16546 50924
rect 56410 50912 56416 50924
rect 16540 50884 56416 50912
rect 16540 50872 16546 50884
rect 56410 50872 56416 50884
rect 56468 50872 56474 50924
rect 57238 50872 57244 50924
rect 57296 50912 57302 50924
rect 64846 50912 64874 50952
rect 78766 50940 78772 50952
rect 78824 50940 78830 50992
rect 81342 50940 81348 50992
rect 81400 50980 81406 50992
rect 85577 50983 85635 50989
rect 85577 50980 85589 50983
rect 81400 50952 85589 50980
rect 81400 50940 81406 50952
rect 85577 50949 85589 50952
rect 85623 50949 85635 50983
rect 85776 50980 85804 51088
rect 85853 51051 85911 51057
rect 85853 51017 85865 51051
rect 85899 51048 85911 51051
rect 112254 51048 112260 51060
rect 85899 51020 112260 51048
rect 85899 51017 85911 51020
rect 85853 51011 85911 51017
rect 112254 51008 112260 51020
rect 112312 51008 112318 51060
rect 115842 51008 115848 51060
rect 115900 51048 115906 51060
rect 141786 51048 141792 51060
rect 115900 51020 141792 51048
rect 115900 51008 115906 51020
rect 141786 51008 141792 51020
rect 141844 51008 141850 51060
rect 144638 51008 144644 51060
rect 144696 51048 144702 51060
rect 166166 51048 166172 51060
rect 144696 51020 166172 51048
rect 144696 51008 144702 51020
rect 166166 51008 166172 51020
rect 166224 51008 166230 51060
rect 168282 51008 168288 51060
rect 168340 51048 168346 51060
rect 186498 51048 186504 51060
rect 168340 51020 186504 51048
rect 168340 51008 168346 51020
rect 186498 51008 186504 51020
rect 186556 51008 186562 51060
rect 190362 51008 190368 51060
rect 190420 51048 190426 51060
rect 205726 51048 205732 51060
rect 190420 51020 205732 51048
rect 190420 51008 190426 51020
rect 205726 51008 205732 51020
rect 205784 51008 205790 51060
rect 208302 51008 208308 51060
rect 208360 51048 208366 51060
rect 220998 51048 221004 51060
rect 208360 51020 221004 51048
rect 208360 51008 208366 51020
rect 220998 51008 221004 51020
rect 221056 51008 221062 51060
rect 222102 51008 222108 51060
rect 222160 51048 222166 51060
rect 233142 51048 233148 51060
rect 222160 51020 233148 51048
rect 222160 51008 222166 51020
rect 233142 51008 233148 51020
rect 233200 51008 233206 51060
rect 530854 51008 530860 51060
rect 530912 51048 530918 51060
rect 544378 51048 544384 51060
rect 530912 51020 544384 51048
rect 530912 51008 530918 51020
rect 544378 51008 544384 51020
rect 544436 51008 544442 51060
rect 109218 50980 109224 50992
rect 85776 50952 109224 50980
rect 85577 50943 85635 50949
rect 109218 50940 109224 50952
rect 109276 50940 109282 50992
rect 113082 50940 113088 50992
rect 113140 50980 113146 50992
rect 139762 50980 139768 50992
rect 113140 50952 139768 50980
rect 113140 50940 113146 50952
rect 139762 50940 139768 50952
rect 139820 50940 139826 50992
rect 140682 50940 140688 50992
rect 140740 50980 140746 50992
rect 163130 50980 163136 50992
rect 140740 50952 163136 50980
rect 140740 50940 140746 50952
rect 163130 50940 163136 50952
rect 163188 50940 163194 50992
rect 166077 50983 166135 50989
rect 166077 50949 166089 50983
rect 166123 50980 166135 50983
rect 173161 50983 173219 50989
rect 173161 50980 173173 50983
rect 166123 50952 173173 50980
rect 166123 50949 166135 50952
rect 166077 50943 166135 50949
rect 173161 50949 173173 50952
rect 173207 50949 173219 50983
rect 173161 50943 173219 50949
rect 173253 50983 173311 50989
rect 173253 50949 173265 50983
rect 173299 50980 173311 50983
rect 182358 50980 182364 50992
rect 173299 50952 182364 50980
rect 173299 50949 173311 50952
rect 173253 50943 173311 50949
rect 182358 50940 182364 50952
rect 182416 50940 182422 50992
rect 183462 50940 183468 50992
rect 183520 50980 183526 50992
rect 199654 50980 199660 50992
rect 183520 50952 199660 50980
rect 183520 50940 183526 50952
rect 199654 50940 199660 50952
rect 199712 50940 199718 50992
rect 200022 50940 200028 50992
rect 200080 50980 200086 50992
rect 213914 50980 213920 50992
rect 200080 50952 213920 50980
rect 200080 50940 200086 50952
rect 213914 50940 213920 50952
rect 213972 50940 213978 50992
rect 215202 50940 215208 50992
rect 215260 50980 215266 50992
rect 227070 50980 227076 50992
rect 215260 50952 227076 50980
rect 215260 50940 215266 50952
rect 227070 50940 227076 50952
rect 227128 50940 227134 50992
rect 227622 50940 227628 50992
rect 227680 50980 227686 50992
rect 237282 50980 237288 50992
rect 227680 50952 237288 50980
rect 227680 50940 227686 50952
rect 237282 50940 237288 50952
rect 237340 50940 237346 50992
rect 241422 50940 241428 50992
rect 241480 50980 241486 50992
rect 249426 50980 249432 50992
rect 241480 50952 249432 50980
rect 241480 50940 241486 50952
rect 249426 50940 249432 50952
rect 249484 50940 249490 50992
rect 252370 50940 252376 50992
rect 252428 50980 252434 50992
rect 259638 50980 259644 50992
rect 252428 50952 259644 50980
rect 252428 50940 252434 50952
rect 259638 50940 259644 50952
rect 259696 50940 259702 50992
rect 510522 50940 510528 50992
rect 510580 50980 510586 50992
rect 536098 50980 536104 50992
rect 510580 50952 536104 50980
rect 510580 50940 510586 50952
rect 536098 50940 536104 50952
rect 536156 50940 536162 50992
rect 57296 50884 64874 50912
rect 57296 50872 57302 50884
rect 67542 50872 67548 50924
rect 67600 50912 67606 50924
rect 67600 50884 68232 50912
rect 67600 50872 67606 50884
rect 12342 50804 12348 50856
rect 12400 50844 12406 50856
rect 52362 50844 52368 50856
rect 12400 50816 52368 50844
rect 12400 50804 12406 50816
rect 52362 50804 52368 50816
rect 52420 50804 52426 50856
rect 56502 50804 56508 50856
rect 56560 50844 56566 50856
rect 63681 50847 63739 50853
rect 63681 50844 63693 50847
rect 56560 50816 63693 50844
rect 56560 50804 56566 50816
rect 63681 50813 63693 50816
rect 63727 50813 63739 50847
rect 63681 50807 63739 50813
rect 63773 50847 63831 50853
rect 63773 50813 63785 50847
rect 63819 50844 63831 50847
rect 67634 50844 67640 50856
rect 63819 50816 67640 50844
rect 63819 50813 63831 50816
rect 63773 50807 63831 50813
rect 67634 50804 67640 50816
rect 67692 50804 67698 50856
rect 20622 50736 20628 50788
rect 20680 50776 20686 50788
rect 59446 50776 59452 50788
rect 20680 50748 59452 50776
rect 20680 50736 20686 50748
rect 59446 50736 59452 50748
rect 59504 50736 59510 50788
rect 63402 50736 63408 50788
rect 63460 50776 63466 50788
rect 68204 50776 68232 50884
rect 70302 50872 70308 50924
rect 70360 50912 70366 50924
rect 103146 50912 103152 50924
rect 70360 50884 103152 50912
rect 70360 50872 70366 50884
rect 103146 50872 103152 50884
rect 103204 50872 103210 50924
rect 110322 50872 110328 50924
rect 110380 50912 110386 50924
rect 136634 50912 136640 50924
rect 110380 50884 136640 50912
rect 110380 50872 110386 50884
rect 136634 50872 136640 50884
rect 136692 50872 136698 50924
rect 139302 50872 139308 50924
rect 139360 50912 139366 50924
rect 162026 50912 162032 50924
rect 139360 50884 162032 50912
rect 139360 50872 139366 50884
rect 162026 50872 162032 50884
rect 162084 50872 162090 50924
rect 165522 50872 165528 50924
rect 165580 50912 165586 50924
rect 184382 50912 184388 50924
rect 165580 50884 184388 50912
rect 165580 50872 165586 50884
rect 184382 50872 184388 50884
rect 184440 50872 184446 50924
rect 186222 50872 186228 50924
rect 186280 50912 186286 50924
rect 201678 50912 201684 50924
rect 186280 50884 201684 50912
rect 186280 50872 186286 50884
rect 201678 50872 201684 50884
rect 201736 50872 201742 50924
rect 205542 50872 205548 50924
rect 205600 50912 205606 50924
rect 218974 50912 218980 50924
rect 205600 50884 218980 50912
rect 205600 50872 205606 50884
rect 218974 50872 218980 50884
rect 219032 50872 219038 50924
rect 219250 50872 219256 50924
rect 219308 50912 219314 50924
rect 230106 50912 230112 50924
rect 219308 50884 230112 50912
rect 219308 50872 219314 50884
rect 230106 50872 230112 50884
rect 230164 50872 230170 50924
rect 234522 50872 234528 50924
rect 234580 50912 234586 50924
rect 243354 50912 243360 50924
rect 234580 50884 243360 50912
rect 234580 50872 234586 50884
rect 243354 50872 243360 50884
rect 243412 50872 243418 50924
rect 253842 50872 253848 50924
rect 253900 50912 253906 50924
rect 260650 50912 260656 50924
rect 253900 50884 260656 50912
rect 253900 50872 253906 50884
rect 260650 50872 260656 50884
rect 260708 50872 260714 50924
rect 509510 50872 509516 50924
rect 509568 50912 509574 50924
rect 542354 50912 542360 50924
rect 509568 50884 542360 50912
rect 509568 50872 509574 50884
rect 542354 50872 542360 50884
rect 542412 50872 542418 50924
rect 68922 50804 68928 50856
rect 68980 50844 68986 50856
rect 101122 50844 101128 50856
rect 68980 50816 101128 50844
rect 68980 50804 68986 50816
rect 101122 50804 101128 50816
rect 101180 50804 101186 50856
rect 107562 50804 107568 50856
rect 107620 50844 107626 50856
rect 134610 50844 134616 50856
rect 107620 50816 134616 50844
rect 107620 50804 107626 50816
rect 134610 50804 134616 50816
rect 134668 50804 134674 50856
rect 144730 50804 144736 50856
rect 144788 50844 144794 50856
rect 167178 50844 167184 50856
rect 144788 50816 167184 50844
rect 144788 50804 144794 50816
rect 167178 50804 167184 50816
rect 167236 50804 167242 50856
rect 173161 50847 173219 50853
rect 173161 50813 173173 50847
rect 173207 50844 173219 50847
rect 179322 50844 179328 50856
rect 173207 50816 179328 50844
rect 173207 50813 173219 50816
rect 173161 50807 173219 50813
rect 179322 50804 179328 50816
rect 179380 50804 179386 50856
rect 180058 50804 180064 50856
rect 180116 50844 180122 50856
rect 180521 50847 180579 50853
rect 180116 50816 180472 50844
rect 180116 50804 180122 50816
rect 100110 50776 100116 50788
rect 63460 50748 68140 50776
rect 68204 50748 100116 50776
rect 63460 50736 63466 50748
rect 10962 50668 10968 50720
rect 11020 50708 11026 50720
rect 51350 50708 51356 50720
rect 11020 50680 51356 50708
rect 11020 50668 11026 50680
rect 51350 50668 51356 50680
rect 51408 50668 51414 50720
rect 54478 50668 54484 50720
rect 54536 50708 54542 50720
rect 63494 50708 63500 50720
rect 54536 50680 63500 50708
rect 54536 50668 54542 50680
rect 63494 50668 63500 50680
rect 63552 50668 63558 50720
rect 67913 50711 67971 50717
rect 67913 50708 67925 50711
rect 63604 50680 67925 50708
rect 15102 50600 15108 50652
rect 15160 50640 15166 50652
rect 55398 50640 55404 50652
rect 15160 50612 55404 50640
rect 15160 50600 15166 50612
rect 55398 50600 55404 50612
rect 55456 50600 55462 50652
rect 55858 50600 55864 50652
rect 55916 50640 55922 50652
rect 58529 50643 58587 50649
rect 58529 50640 58541 50643
rect 55916 50612 58541 50640
rect 55916 50600 55922 50612
rect 58529 50609 58541 50612
rect 58575 50609 58587 50643
rect 58529 50603 58587 50609
rect 13722 50532 13728 50584
rect 13780 50572 13786 50584
rect 54386 50572 54392 50584
rect 13780 50544 54392 50572
rect 13780 50532 13786 50544
rect 54386 50532 54392 50544
rect 54444 50532 54450 50584
rect 60642 50532 60648 50584
rect 60700 50572 60706 50584
rect 63604 50572 63632 50680
rect 67913 50677 67925 50680
rect 67959 50677 67971 50711
rect 67913 50671 67971 50677
rect 63773 50643 63831 50649
rect 63773 50609 63785 50643
rect 63819 50640 63831 50643
rect 66530 50640 66536 50652
rect 63819 50612 66536 50640
rect 63819 50609 63831 50612
rect 63773 50603 63831 50609
rect 66530 50600 66536 50612
rect 66588 50600 66594 50652
rect 68112 50640 68140 50748
rect 100110 50736 100116 50748
rect 100168 50736 100174 50788
rect 103422 50736 103428 50788
rect 103480 50776 103486 50788
rect 130562 50776 130568 50788
rect 103480 50748 130568 50776
rect 103480 50736 103486 50748
rect 130562 50736 130568 50748
rect 130620 50736 130626 50788
rect 137922 50736 137928 50788
rect 137980 50776 137986 50788
rect 161014 50776 161020 50788
rect 137980 50748 161020 50776
rect 137980 50736 137986 50748
rect 161014 50736 161020 50748
rect 161072 50736 161078 50788
rect 161382 50736 161388 50788
rect 161440 50776 161446 50788
rect 166169 50779 166227 50785
rect 166169 50776 166181 50779
rect 161440 50748 166181 50776
rect 161440 50736 161446 50748
rect 166169 50745 166181 50748
rect 166215 50745 166227 50779
rect 166169 50739 166227 50745
rect 166353 50779 166411 50785
rect 166353 50745 166365 50779
rect 166399 50776 166411 50779
rect 180334 50776 180340 50788
rect 166399 50748 180340 50776
rect 166399 50745 166411 50748
rect 166353 50739 166411 50745
rect 180334 50736 180340 50748
rect 180392 50736 180398 50788
rect 180444 50776 180472 50816
rect 180521 50813 180533 50847
rect 180567 50844 180579 50847
rect 190546 50844 190552 50856
rect 180567 50816 190552 50844
rect 180567 50813 180579 50816
rect 180521 50807 180579 50813
rect 190546 50804 190552 50816
rect 190604 50804 190610 50856
rect 194410 50804 194416 50856
rect 194468 50844 194474 50856
rect 208762 50844 208768 50856
rect 194468 50816 208768 50844
rect 194468 50804 194474 50816
rect 208762 50804 208768 50816
rect 208820 50804 208826 50856
rect 211062 50804 211068 50856
rect 211120 50844 211126 50856
rect 223022 50844 223028 50856
rect 211120 50816 223028 50844
rect 211120 50804 211126 50816
rect 223022 50804 223028 50816
rect 223080 50804 223086 50856
rect 223482 50804 223488 50856
rect 223540 50844 223546 50856
rect 234246 50844 234252 50856
rect 223540 50816 234252 50844
rect 223540 50804 223546 50816
rect 234246 50804 234252 50816
rect 234304 50804 234310 50856
rect 235902 50804 235908 50856
rect 235960 50844 235966 50856
rect 244366 50844 244372 50856
rect 235960 50816 244372 50844
rect 235960 50804 235966 50816
rect 244366 50804 244372 50816
rect 244424 50804 244430 50856
rect 262122 50804 262128 50856
rect 262180 50844 262186 50856
rect 267734 50844 267740 50856
rect 262180 50816 267740 50844
rect 262180 50804 262186 50816
rect 267734 50804 267740 50816
rect 267792 50804 267798 50856
rect 506474 50804 506480 50856
rect 506532 50844 506538 50856
rect 533341 50847 533399 50853
rect 533341 50844 533353 50847
rect 506532 50816 533353 50844
rect 506532 50804 506538 50816
rect 533341 50813 533353 50816
rect 533387 50813 533399 50847
rect 533341 50807 533399 50813
rect 542998 50804 543004 50856
rect 543056 50844 543062 50856
rect 548518 50844 548524 50856
rect 543056 50816 548524 50844
rect 543056 50804 543062 50816
rect 548518 50804 548524 50816
rect 548576 50804 548582 50856
rect 181346 50776 181352 50788
rect 180444 50748 181352 50776
rect 181346 50736 181352 50748
rect 181404 50736 181410 50788
rect 197630 50776 197636 50788
rect 185596 50748 197636 50776
rect 68189 50711 68247 50717
rect 68189 50677 68201 50711
rect 68235 50708 68247 50711
rect 88981 50711 89039 50717
rect 88981 50708 88993 50711
rect 68235 50680 88993 50708
rect 68235 50677 68247 50680
rect 68189 50671 68247 50677
rect 88981 50677 88993 50680
rect 89027 50677 89039 50711
rect 88981 50671 89039 50677
rect 89070 50668 89076 50720
rect 89128 50708 89134 50720
rect 95050 50708 95056 50720
rect 89128 50680 95056 50708
rect 89128 50668 89134 50680
rect 95050 50668 95056 50680
rect 95108 50668 95114 50720
rect 95142 50668 95148 50720
rect 95200 50708 95206 50720
rect 97813 50711 97871 50717
rect 97813 50708 97825 50711
rect 95200 50680 97825 50708
rect 95200 50668 95206 50680
rect 97813 50677 97825 50680
rect 97859 50677 97871 50711
rect 97813 50671 97871 50677
rect 99282 50668 99288 50720
rect 99340 50708 99346 50720
rect 127526 50708 127532 50720
rect 99340 50680 127532 50708
rect 99340 50668 99346 50680
rect 127526 50668 127532 50680
rect 127584 50668 127590 50720
rect 136542 50668 136548 50720
rect 136600 50708 136606 50720
rect 158990 50708 158996 50720
rect 136600 50680 158996 50708
rect 136600 50668 136606 50680
rect 158990 50668 158996 50680
rect 159048 50668 159054 50720
rect 160002 50668 160008 50720
rect 160060 50708 160066 50720
rect 166077 50711 166135 50717
rect 166077 50708 166089 50711
rect 160060 50680 166089 50708
rect 160060 50668 160066 50680
rect 166077 50677 166089 50680
rect 166123 50677 166135 50711
rect 166077 50671 166135 50677
rect 166902 50668 166908 50720
rect 166960 50708 166966 50720
rect 185394 50708 185400 50720
rect 166960 50680 185400 50708
rect 166960 50668 166966 50680
rect 185394 50668 185400 50680
rect 185452 50668 185458 50720
rect 97074 50640 97080 50652
rect 68112 50612 97080 50640
rect 97074 50600 97080 50612
rect 97132 50600 97138 50652
rect 100662 50600 100668 50652
rect 100720 50640 100726 50652
rect 128538 50640 128544 50652
rect 100720 50612 128544 50640
rect 100720 50600 100726 50612
rect 128538 50600 128544 50612
rect 128596 50600 128602 50652
rect 135162 50600 135168 50652
rect 135220 50640 135226 50652
rect 157978 50640 157984 50652
rect 135220 50612 157984 50640
rect 135220 50600 135226 50612
rect 157978 50600 157984 50612
rect 158036 50600 158042 50652
rect 162762 50600 162768 50652
rect 162820 50640 162826 50652
rect 173253 50643 173311 50649
rect 173253 50640 173265 50643
rect 162820 50612 173265 50640
rect 162820 50600 162826 50612
rect 173253 50609 173265 50612
rect 173299 50609 173311 50643
rect 173253 50603 173311 50609
rect 180702 50600 180708 50652
rect 180760 50640 180766 50652
rect 185596 50640 185624 50748
rect 197630 50736 197636 50748
rect 197688 50736 197694 50788
rect 198642 50736 198648 50788
rect 198700 50776 198706 50788
rect 212902 50776 212908 50788
rect 198700 50748 212908 50776
rect 198700 50736 198706 50748
rect 212902 50736 212908 50748
rect 212960 50736 212966 50788
rect 213822 50736 213828 50788
rect 213880 50776 213886 50788
rect 226058 50776 226064 50788
rect 213880 50748 226064 50776
rect 213880 50736 213886 50748
rect 226058 50736 226064 50748
rect 226116 50736 226122 50788
rect 226242 50736 226248 50788
rect 226300 50776 226306 50788
rect 236270 50776 236276 50788
rect 226300 50748 236276 50776
rect 226300 50736 226306 50748
rect 236270 50736 236276 50748
rect 236328 50736 236334 50788
rect 237282 50736 237288 50788
rect 237340 50776 237346 50788
rect 246390 50776 246396 50788
rect 237340 50748 246396 50776
rect 237340 50736 237346 50748
rect 246390 50736 246396 50748
rect 246448 50736 246454 50788
rect 246942 50736 246948 50788
rect 247000 50776 247006 50788
rect 254486 50776 254492 50788
rect 247000 50748 254492 50776
rect 247000 50736 247006 50748
rect 254486 50736 254492 50748
rect 254544 50736 254550 50788
rect 264882 50736 264888 50788
rect 264940 50776 264946 50788
rect 269758 50776 269764 50788
rect 264940 50748 269764 50776
rect 264940 50736 264946 50748
rect 269758 50736 269764 50748
rect 269816 50736 269822 50788
rect 275922 50736 275928 50788
rect 275980 50776 275986 50788
rect 278866 50776 278872 50788
rect 275980 50748 278872 50776
rect 275980 50736 275986 50748
rect 278866 50736 278872 50748
rect 278924 50736 278930 50788
rect 285490 50736 285496 50788
rect 285548 50776 285554 50788
rect 288066 50776 288072 50788
rect 285548 50748 288072 50776
rect 285548 50736 285554 50748
rect 288066 50736 288072 50748
rect 288124 50736 288130 50788
rect 332778 50736 332784 50788
rect 332836 50776 332842 50788
rect 335998 50776 336004 50788
rect 332836 50748 336004 50776
rect 332836 50736 332842 50748
rect 335998 50736 336004 50748
rect 336056 50736 336062 50788
rect 458726 50736 458732 50788
rect 458784 50776 458790 50788
rect 461578 50776 461584 50788
rect 458784 50748 461584 50776
rect 458784 50736 458790 50748
rect 461578 50736 461584 50748
rect 461636 50736 461642 50788
rect 477034 50736 477040 50788
rect 477092 50776 477098 50788
rect 482278 50776 482284 50788
rect 477092 50748 482284 50776
rect 477092 50736 477098 50748
rect 482278 50736 482284 50748
rect 482336 50736 482342 50788
rect 516594 50736 516600 50788
rect 516652 50776 516658 50788
rect 520918 50776 520924 50788
rect 516652 50748 520924 50776
rect 516652 50736 516658 50748
rect 520918 50736 520924 50748
rect 520976 50736 520982 50788
rect 522758 50736 522764 50788
rect 522816 50776 522822 50788
rect 556798 50776 556804 50788
rect 522816 50748 556804 50776
rect 522816 50736 522822 50748
rect 556798 50736 556804 50748
rect 556856 50736 556862 50788
rect 187602 50668 187608 50720
rect 187660 50708 187666 50720
rect 203702 50708 203708 50720
rect 187660 50680 203708 50708
rect 187660 50668 187666 50680
rect 203702 50668 203708 50680
rect 203760 50668 203766 50720
rect 204162 50668 204168 50720
rect 204220 50708 204226 50720
rect 217962 50708 217968 50720
rect 204220 50680 217968 50708
rect 204220 50668 204226 50680
rect 217962 50668 217968 50680
rect 218020 50668 218026 50720
rect 219342 50668 219348 50720
rect 219400 50708 219406 50720
rect 231118 50708 231124 50720
rect 219400 50680 231124 50708
rect 219400 50668 219406 50680
rect 231118 50668 231124 50680
rect 231176 50668 231182 50720
rect 231762 50668 231768 50720
rect 231820 50708 231826 50720
rect 241330 50708 241336 50720
rect 231820 50680 241336 50708
rect 231820 50668 231826 50680
rect 241330 50668 241336 50680
rect 241388 50668 241394 50720
rect 244182 50668 244188 50720
rect 244240 50708 244246 50720
rect 252462 50708 252468 50720
rect 244240 50680 252468 50708
rect 244240 50668 244246 50680
rect 252462 50668 252468 50680
rect 252520 50668 252526 50720
rect 267642 50668 267648 50720
rect 267700 50708 267706 50720
rect 271782 50708 271788 50720
rect 267700 50680 271788 50708
rect 267700 50668 267706 50680
rect 271782 50668 271788 50680
rect 271840 50668 271846 50720
rect 277302 50668 277308 50720
rect 277360 50708 277366 50720
rect 279878 50708 279884 50720
rect 277360 50680 279884 50708
rect 277360 50668 277366 50680
rect 279878 50668 279884 50680
rect 279936 50668 279942 50720
rect 285582 50668 285588 50720
rect 285640 50708 285646 50720
rect 287054 50708 287060 50720
rect 285640 50680 287060 50708
rect 285640 50668 285646 50680
rect 287054 50668 287060 50680
rect 287112 50668 287118 50720
rect 525794 50668 525800 50720
rect 525852 50708 525858 50720
rect 560938 50708 560944 50720
rect 525852 50680 560944 50708
rect 525852 50668 525858 50680
rect 560938 50668 560944 50680
rect 560996 50668 561002 50720
rect 180760 50612 185624 50640
rect 180760 50600 180766 50612
rect 186130 50600 186136 50652
rect 186188 50640 186194 50652
rect 202690 50640 202696 50652
rect 186188 50612 202696 50640
rect 186188 50600 186194 50612
rect 202690 50600 202696 50612
rect 202748 50600 202754 50652
rect 202782 50600 202788 50652
rect 202840 50640 202846 50652
rect 215938 50640 215944 50652
rect 202840 50612 215944 50640
rect 202840 50600 202846 50612
rect 215938 50600 215944 50612
rect 215996 50600 216002 50652
rect 216582 50600 216588 50652
rect 216640 50640 216646 50652
rect 228082 50640 228088 50652
rect 216640 50612 228088 50640
rect 216640 50600 216646 50612
rect 228082 50600 228088 50612
rect 228140 50600 228146 50652
rect 229002 50600 229008 50652
rect 229060 50640 229066 50652
rect 239306 50640 239312 50652
rect 229060 50612 239312 50640
rect 229060 50600 229066 50612
rect 239306 50600 239312 50612
rect 239364 50600 239370 50652
rect 240042 50600 240048 50652
rect 240100 50640 240106 50652
rect 248414 50640 248420 50652
rect 240100 50612 248420 50640
rect 240100 50600 240106 50612
rect 248414 50600 248420 50612
rect 248472 50600 248478 50652
rect 256602 50600 256608 50652
rect 256660 50640 256666 50652
rect 262674 50640 262680 50652
rect 256660 50612 262680 50640
rect 256660 50600 256666 50612
rect 262674 50600 262680 50612
rect 262732 50600 262738 50652
rect 274542 50600 274548 50652
rect 274600 50640 274606 50652
rect 277854 50640 277860 50652
rect 274600 50612 277860 50640
rect 274600 50600 274606 50612
rect 277854 50600 277860 50612
rect 277912 50600 277918 50652
rect 492214 50600 492220 50652
rect 492272 50640 492278 50652
rect 500218 50640 500224 50652
rect 492272 50612 500224 50640
rect 492272 50600 492278 50612
rect 500218 50600 500224 50612
rect 500276 50600 500282 50652
rect 528830 50600 528836 50652
rect 528888 50640 528894 50652
rect 564526 50640 564532 50652
rect 528888 50612 564532 50640
rect 528888 50600 528894 50612
rect 564526 50600 564532 50612
rect 564584 50600 564590 50652
rect 60700 50544 63632 50572
rect 63681 50575 63739 50581
rect 60700 50532 60706 50544
rect 63681 50541 63693 50575
rect 63727 50572 63739 50575
rect 91002 50572 91008 50584
rect 63727 50544 91008 50572
rect 63727 50541 63739 50544
rect 63681 50535 63739 50541
rect 91002 50532 91008 50544
rect 91060 50532 91066 50584
rect 119430 50572 119436 50584
rect 91204 50544 119436 50572
rect 9582 50464 9588 50516
rect 9640 50504 9646 50516
rect 50338 50504 50344 50516
rect 9640 50476 50344 50504
rect 9640 50464 9646 50476
rect 50338 50464 50344 50476
rect 50396 50464 50402 50516
rect 53742 50464 53748 50516
rect 53800 50504 53806 50516
rect 87874 50504 87880 50516
rect 53800 50476 87880 50504
rect 53800 50464 53806 50476
rect 87874 50464 87880 50476
rect 87932 50464 87938 50516
rect 88981 50507 89039 50513
rect 88981 50473 88993 50507
rect 89027 50504 89039 50507
rect 91097 50507 91155 50513
rect 91097 50504 91109 50507
rect 89027 50476 91109 50504
rect 89027 50473 89039 50476
rect 88981 50467 89039 50473
rect 91097 50473 91109 50476
rect 91143 50473 91155 50507
rect 91097 50467 91155 50473
rect 6822 50396 6828 50448
rect 6880 50436 6886 50448
rect 48314 50436 48320 50448
rect 6880 50408 48320 50436
rect 6880 50396 6886 50408
rect 48314 50396 48320 50408
rect 48372 50396 48378 50448
rect 50982 50396 50988 50448
rect 51040 50436 51046 50448
rect 85850 50436 85856 50448
rect 51040 50408 85856 50436
rect 51040 50396 51046 50408
rect 85850 50396 85856 50408
rect 85908 50396 85914 50448
rect 90358 50396 90364 50448
rect 90416 50436 90422 50448
rect 91204 50436 91232 50544
rect 119430 50532 119436 50544
rect 119488 50532 119494 50584
rect 119982 50532 119988 50584
rect 120040 50572 120046 50584
rect 145834 50572 145840 50584
rect 120040 50544 145840 50572
rect 120040 50532 120046 50544
rect 145834 50532 145840 50544
rect 145892 50532 145898 50584
rect 146938 50532 146944 50584
rect 146996 50572 147002 50584
rect 152918 50572 152924 50584
rect 146996 50544 152924 50572
rect 146996 50532 147002 50544
rect 152918 50532 152924 50544
rect 152976 50532 152982 50584
rect 153013 50575 153071 50581
rect 153013 50541 153025 50575
rect 153059 50572 153071 50575
rect 168190 50572 168196 50584
rect 153059 50544 168196 50572
rect 153059 50541 153071 50544
rect 153013 50535 153071 50541
rect 168190 50532 168196 50544
rect 168248 50532 168254 50584
rect 169662 50532 169668 50584
rect 169720 50572 169726 50584
rect 188522 50572 188528 50584
rect 169720 50544 188528 50572
rect 169720 50532 169726 50544
rect 188522 50532 188528 50544
rect 188580 50532 188586 50584
rect 188982 50532 188988 50584
rect 189040 50572 189046 50584
rect 204714 50572 204720 50584
rect 189040 50544 204720 50572
rect 189040 50532 189046 50544
rect 204714 50532 204720 50544
rect 204772 50532 204778 50584
rect 206922 50532 206928 50584
rect 206980 50572 206986 50584
rect 219986 50572 219992 50584
rect 206980 50544 219992 50572
rect 206980 50532 206986 50544
rect 219986 50532 219992 50544
rect 220044 50532 220050 50584
rect 220722 50532 220728 50584
rect 220780 50572 220786 50584
rect 232130 50572 232136 50584
rect 220780 50544 232136 50572
rect 220780 50532 220786 50544
rect 232130 50532 232136 50544
rect 232188 50532 232194 50584
rect 233142 50532 233148 50584
rect 233200 50572 233206 50584
rect 242342 50572 242348 50584
rect 233200 50544 242348 50572
rect 233200 50532 233206 50544
rect 242342 50532 242348 50544
rect 242400 50532 242406 50584
rect 242802 50532 242808 50584
rect 242860 50572 242866 50584
rect 250438 50572 250444 50584
rect 242860 50544 250444 50572
rect 242860 50532 242866 50544
rect 250438 50532 250444 50544
rect 250496 50532 250502 50584
rect 266998 50532 267004 50584
rect 267056 50572 267062 50584
rect 270770 50572 270776 50584
rect 267056 50544 270776 50572
rect 267056 50532 267062 50544
rect 270770 50532 270776 50544
rect 270828 50532 270834 50584
rect 286962 50532 286968 50584
rect 287020 50572 287026 50584
rect 289078 50572 289084 50584
rect 287020 50544 289084 50572
rect 287020 50532 287026 50544
rect 289078 50532 289084 50544
rect 289136 50532 289142 50584
rect 495250 50532 495256 50584
rect 495308 50572 495314 50584
rect 504358 50572 504364 50584
rect 495308 50544 504364 50572
rect 495308 50532 495314 50544
rect 504358 50532 504364 50544
rect 504416 50532 504422 50584
rect 519630 50532 519636 50584
rect 519688 50572 519694 50584
rect 554774 50572 554780 50584
rect 519688 50544 554780 50572
rect 519688 50532 519694 50544
rect 554774 50532 554780 50544
rect 554832 50532 554838 50584
rect 91281 50507 91339 50513
rect 91281 50473 91293 50507
rect 91327 50504 91339 50507
rect 94038 50504 94044 50516
rect 91327 50476 94044 50504
rect 91327 50473 91339 50476
rect 91281 50467 91339 50473
rect 94038 50464 94044 50476
rect 94096 50464 94102 50516
rect 97721 50507 97779 50513
rect 97721 50473 97733 50507
rect 97767 50504 97779 50507
rect 118418 50504 118424 50516
rect 97767 50476 118424 50504
rect 97767 50473 97779 50476
rect 97721 50467 97779 50473
rect 118418 50464 118424 50476
rect 118476 50464 118482 50516
rect 121362 50464 121368 50516
rect 121420 50504 121426 50516
rect 146846 50504 146852 50516
rect 121420 50476 146852 50504
rect 121420 50464 121426 50476
rect 146846 50464 146852 50476
rect 146904 50464 146910 50516
rect 148962 50464 148968 50516
rect 149020 50504 149026 50516
rect 170214 50504 170220 50516
rect 149020 50476 170220 50504
rect 149020 50464 149026 50476
rect 170214 50464 170220 50476
rect 170272 50464 170278 50516
rect 171042 50464 171048 50516
rect 171100 50504 171106 50516
rect 189534 50504 189540 50516
rect 171100 50476 189540 50504
rect 171100 50464 171106 50476
rect 189534 50464 189540 50476
rect 189592 50464 189598 50516
rect 194502 50464 194508 50516
rect 194560 50504 194566 50516
rect 209774 50504 209780 50516
rect 194560 50476 209780 50504
rect 194560 50464 194566 50476
rect 209774 50464 209780 50476
rect 209832 50464 209838 50516
rect 210970 50464 210976 50516
rect 211028 50504 211034 50516
rect 224034 50504 224040 50516
rect 211028 50476 224040 50504
rect 211028 50464 211034 50476
rect 224034 50464 224040 50476
rect 224092 50464 224098 50516
rect 224862 50464 224868 50516
rect 224920 50504 224926 50516
rect 235258 50504 235264 50516
rect 224920 50476 235264 50504
rect 224920 50464 224926 50476
rect 235258 50464 235264 50476
rect 235316 50464 235322 50516
rect 235810 50464 235816 50516
rect 235868 50504 235874 50516
rect 245378 50504 245384 50516
rect 235868 50476 245384 50504
rect 235868 50464 235874 50476
rect 245378 50464 245384 50476
rect 245436 50464 245442 50516
rect 245562 50464 245568 50516
rect 245620 50504 245626 50516
rect 253474 50504 253480 50516
rect 245620 50476 253480 50504
rect 245620 50464 245626 50476
rect 253474 50464 253480 50476
rect 253532 50464 253538 50516
rect 255222 50464 255228 50516
rect 255280 50504 255286 50516
rect 261662 50504 261668 50516
rect 255280 50476 261668 50504
rect 255280 50464 255286 50476
rect 261662 50464 261668 50476
rect 261720 50464 261726 50516
rect 494238 50464 494244 50516
rect 494296 50504 494302 50516
rect 515398 50504 515404 50516
rect 494296 50476 515404 50504
rect 494296 50464 494302 50476
rect 515398 50464 515404 50476
rect 515456 50464 515462 50516
rect 533341 50507 533399 50513
rect 533341 50473 533353 50507
rect 533387 50504 533399 50507
rect 539594 50504 539600 50516
rect 533387 50476 539600 50504
rect 533387 50473 533399 50476
rect 533341 50467 533399 50473
rect 539594 50464 539600 50476
rect 539652 50464 539658 50516
rect 543001 50507 543059 50513
rect 543001 50473 543013 50507
rect 543047 50504 543059 50507
rect 568574 50504 568580 50516
rect 543047 50476 568580 50504
rect 543047 50473 543059 50476
rect 543001 50467 543059 50473
rect 568574 50464 568580 50476
rect 568632 50464 568638 50516
rect 90416 50408 91232 50436
rect 90416 50396 90422 50408
rect 92382 50396 92388 50448
rect 92440 50436 92446 50448
rect 121454 50436 121460 50448
rect 92440 50408 121460 50436
rect 92440 50396 92446 50408
rect 121454 50396 121460 50408
rect 121512 50396 121518 50448
rect 122742 50396 122748 50448
rect 122800 50436 122806 50448
rect 147858 50436 147864 50448
rect 122800 50408 147864 50436
rect 122800 50396 122806 50408
rect 147858 50396 147864 50408
rect 147916 50396 147922 50448
rect 153010 50396 153016 50448
rect 153068 50436 153074 50448
rect 174262 50436 174268 50448
rect 153068 50408 174268 50436
rect 153068 50396 153074 50408
rect 174262 50396 174268 50408
rect 174320 50396 174326 50448
rect 177850 50396 177856 50448
rect 177908 50436 177914 50448
rect 194594 50436 194600 50448
rect 177908 50408 194600 50436
rect 177908 50396 177914 50408
rect 194594 50396 194600 50408
rect 194652 50396 194658 50448
rect 197262 50396 197268 50448
rect 197320 50436 197326 50448
rect 211890 50436 211896 50448
rect 197320 50408 211896 50436
rect 197320 50396 197326 50408
rect 211890 50396 211896 50408
rect 211948 50396 211954 50448
rect 212442 50396 212448 50448
rect 212500 50436 212506 50448
rect 225046 50436 225052 50448
rect 212500 50408 225052 50436
rect 212500 50396 212506 50408
rect 225046 50396 225052 50408
rect 225104 50396 225110 50448
rect 227530 50396 227536 50448
rect 227588 50436 227594 50448
rect 238294 50436 238300 50448
rect 227588 50408 238300 50436
rect 227588 50396 227594 50408
rect 238294 50396 238300 50408
rect 238352 50396 238358 50448
rect 238662 50396 238668 50448
rect 238720 50436 238726 50448
rect 247402 50436 247408 50448
rect 238720 50408 247408 50436
rect 238720 50396 238726 50408
rect 247402 50396 247408 50408
rect 247460 50396 247466 50448
rect 248322 50396 248328 50448
rect 248380 50436 248386 50448
rect 255498 50436 255504 50448
rect 248380 50408 255504 50436
rect 248380 50396 248386 50408
rect 255498 50396 255504 50408
rect 255556 50396 255562 50448
rect 257982 50396 257988 50448
rect 258040 50436 258046 50448
rect 263686 50436 263692 50448
rect 258040 50408 263692 50436
rect 258040 50396 258046 50408
rect 263686 50396 263692 50408
rect 263744 50396 263750 50448
rect 488166 50396 488172 50448
rect 488224 50436 488230 50448
rect 497458 50436 497464 50448
rect 488224 50408 497464 50436
rect 488224 50396 488230 50408
rect 497458 50396 497464 50408
rect 497516 50396 497522 50448
rect 498378 50396 498384 50448
rect 498436 50436 498442 50448
rect 525058 50436 525064 50448
rect 498436 50408 525064 50436
rect 498436 50396 498442 50408
rect 525058 50396 525064 50408
rect 525116 50396 525122 50448
rect 537938 50396 537944 50448
rect 537996 50436 538002 50448
rect 575474 50436 575480 50448
rect 537996 50408 575480 50436
rect 537996 50396 538002 50408
rect 575474 50396 575480 50408
rect 575532 50396 575538 50448
rect 4062 50328 4068 50380
rect 4120 50368 4126 50380
rect 46290 50368 46296 50380
rect 4120 50340 46296 50368
rect 4120 50328 4126 50340
rect 46290 50328 46296 50340
rect 46348 50328 46354 50380
rect 49602 50328 49608 50380
rect 49660 50368 49666 50380
rect 84838 50368 84844 50380
rect 49660 50340 84844 50368
rect 49660 50328 49666 50340
rect 84838 50328 84844 50340
rect 84896 50328 84902 50380
rect 88242 50328 88248 50380
rect 88300 50368 88306 50380
rect 97721 50371 97779 50377
rect 97721 50368 97733 50371
rect 88300 50340 97733 50368
rect 88300 50328 88306 50340
rect 97721 50337 97733 50340
rect 97767 50337 97779 50371
rect 97721 50331 97779 50337
rect 97813 50371 97871 50377
rect 97813 50337 97825 50371
rect 97859 50368 97871 50371
rect 124490 50368 124496 50380
rect 97859 50340 124496 50368
rect 97859 50337 97871 50340
rect 97813 50331 97871 50337
rect 124490 50328 124496 50340
rect 124548 50328 124554 50380
rect 125413 50371 125471 50377
rect 125413 50337 125425 50371
rect 125459 50368 125471 50371
rect 131574 50368 131580 50380
rect 125459 50340 131580 50368
rect 125459 50337 125471 50340
rect 125413 50331 125471 50337
rect 131574 50328 131580 50340
rect 131632 50328 131638 50380
rect 132402 50328 132408 50380
rect 132460 50368 132466 50380
rect 155954 50368 155960 50380
rect 132460 50340 155960 50368
rect 132460 50328 132466 50340
rect 155954 50328 155960 50340
rect 156012 50328 156018 50380
rect 158622 50328 158628 50380
rect 158680 50368 158686 50380
rect 178310 50368 178316 50380
rect 158680 50340 178316 50368
rect 158680 50328 158686 50340
rect 178310 50328 178316 50340
rect 178368 50328 178374 50380
rect 179322 50328 179328 50380
rect 179380 50368 179386 50380
rect 196618 50368 196624 50380
rect 179380 50340 196624 50368
rect 179380 50328 179386 50340
rect 196618 50328 196624 50340
rect 196676 50328 196682 50380
rect 202782 50328 202788 50380
rect 202840 50368 202846 50380
rect 216950 50368 216956 50380
rect 202840 50340 216956 50368
rect 202840 50328 202846 50340
rect 216950 50328 216956 50340
rect 217008 50328 217014 50380
rect 217962 50328 217968 50380
rect 218020 50368 218026 50380
rect 229094 50368 229100 50380
rect 218020 50340 229100 50368
rect 218020 50328 218026 50340
rect 229094 50328 229100 50340
rect 229152 50328 229158 50380
rect 230382 50328 230388 50380
rect 230440 50368 230446 50380
rect 240318 50368 240324 50380
rect 230440 50340 240324 50368
rect 230440 50328 230446 50340
rect 240318 50328 240324 50340
rect 240376 50328 240382 50380
rect 244090 50328 244096 50380
rect 244148 50368 244154 50380
rect 251450 50368 251456 50380
rect 244148 50340 251456 50368
rect 244148 50328 244154 50340
rect 251450 50328 251456 50340
rect 251508 50328 251514 50380
rect 252462 50328 252468 50380
rect 252520 50368 252526 50380
rect 258626 50368 258632 50380
rect 252520 50340 258632 50368
rect 252520 50328 252526 50340
rect 258626 50328 258632 50340
rect 258684 50328 258690 50380
rect 277210 50328 277216 50380
rect 277268 50368 277274 50380
rect 280890 50368 280896 50380
rect 277268 50340 280896 50368
rect 277268 50328 277274 50340
rect 280890 50328 280896 50340
rect 280948 50328 280954 50380
rect 343910 50328 343916 50380
rect 343968 50368 343974 50380
rect 349246 50368 349252 50380
rect 343968 50340 349252 50368
rect 343968 50328 343974 50340
rect 349246 50328 349252 50340
rect 349304 50328 349310 50380
rect 440418 50328 440424 50380
rect 440476 50368 440482 50380
rect 446398 50368 446404 50380
rect 440476 50340 446404 50368
rect 440476 50328 440482 50340
rect 446398 50328 446404 50340
rect 446456 50328 446462 50380
rect 473998 50328 474004 50380
rect 474056 50368 474062 50380
rect 493318 50368 493324 50380
rect 474056 50340 493324 50368
rect 474056 50328 474062 50340
rect 493318 50328 493324 50340
rect 493376 50328 493382 50380
rect 503438 50328 503444 50380
rect 503496 50368 503502 50380
rect 530578 50368 530584 50380
rect 503496 50340 530584 50368
rect 503496 50328 503502 50340
rect 530578 50328 530584 50340
rect 530636 50328 530642 50380
rect 534902 50328 534908 50380
rect 534960 50368 534966 50380
rect 572806 50368 572812 50380
rect 534960 50340 572812 50368
rect 534960 50328 534966 50340
rect 572806 50328 572812 50340
rect 572864 50328 572870 50380
rect 33042 50260 33048 50312
rect 33100 50300 33106 50312
rect 70670 50300 70676 50312
rect 33100 50272 70676 50300
rect 33100 50260 33106 50272
rect 70670 50260 70676 50272
rect 70728 50260 70734 50312
rect 75822 50260 75828 50312
rect 75880 50300 75886 50312
rect 107194 50300 107200 50312
rect 75880 50272 107200 50300
rect 75880 50260 75886 50272
rect 107194 50260 107200 50272
rect 107252 50260 107258 50312
rect 111702 50260 111708 50312
rect 111760 50300 111766 50312
rect 137646 50300 137652 50312
rect 111760 50272 137652 50300
rect 111760 50260 111766 50272
rect 137646 50260 137652 50272
rect 137704 50260 137710 50312
rect 143442 50260 143448 50312
rect 143500 50300 143506 50312
rect 165154 50300 165160 50312
rect 143500 50272 165160 50300
rect 143500 50260 143506 50272
rect 165154 50260 165160 50272
rect 165212 50260 165218 50312
rect 169570 50260 169576 50312
rect 169628 50300 169634 50312
rect 187510 50300 187516 50312
rect 169628 50272 187516 50300
rect 169628 50260 169634 50272
rect 187510 50260 187516 50272
rect 187568 50260 187574 50312
rect 191742 50260 191748 50312
rect 191800 50300 191806 50312
rect 206738 50300 206744 50312
rect 191800 50272 206744 50300
rect 191800 50260 191806 50272
rect 206738 50260 206744 50272
rect 206796 50260 206802 50312
rect 209682 50260 209688 50312
rect 209740 50300 209746 50312
rect 222010 50300 222016 50312
rect 209740 50272 222016 50300
rect 209740 50260 209746 50272
rect 222010 50260 222016 50272
rect 222068 50260 222074 50312
rect 527818 50260 527824 50312
rect 527876 50300 527882 50312
rect 540238 50300 540244 50312
rect 527876 50272 540244 50300
rect 527876 50260 527882 50272
rect 540238 50260 540244 50272
rect 540296 50260 540302 50312
rect 28902 50192 28908 50244
rect 28960 50232 28966 50244
rect 63773 50235 63831 50241
rect 63773 50232 63785 50235
rect 28960 50204 63785 50232
rect 28960 50192 28966 50204
rect 63773 50201 63785 50204
rect 63819 50201 63831 50235
rect 63773 50195 63831 50201
rect 64138 50192 64144 50244
rect 64196 50232 64202 50244
rect 64196 50204 64874 50232
rect 64196 50192 64202 50204
rect 26142 50124 26148 50176
rect 26200 50164 26206 50176
rect 64506 50164 64512 50176
rect 26200 50136 64512 50164
rect 26200 50124 26206 50136
rect 64506 50124 64512 50136
rect 64564 50124 64570 50176
rect 64846 50164 64874 50204
rect 74442 50192 74448 50244
rect 74500 50232 74506 50244
rect 106182 50232 106188 50244
rect 74500 50204 106188 50232
rect 74500 50192 74506 50204
rect 106182 50192 106188 50204
rect 106240 50192 106246 50244
rect 106274 50192 106280 50244
rect 106332 50232 106338 50244
rect 133598 50232 133604 50244
rect 106332 50204 133604 50232
rect 106332 50192 106338 50204
rect 133598 50192 133604 50204
rect 133656 50192 133662 50244
rect 134518 50192 134524 50244
rect 134576 50232 134582 50244
rect 135622 50232 135628 50244
rect 134576 50204 135628 50232
rect 134576 50192 134582 50204
rect 135622 50192 135628 50204
rect 135680 50192 135686 50244
rect 142062 50192 142068 50244
rect 142120 50232 142126 50244
rect 163774 50232 163780 50244
rect 142120 50204 163780 50232
rect 142120 50192 142126 50204
rect 163774 50192 163780 50204
rect 163832 50192 163838 50244
rect 164142 50192 164148 50244
rect 164200 50232 164206 50244
rect 183370 50232 183376 50244
rect 164200 50204 183376 50232
rect 164200 50192 164206 50204
rect 183370 50192 183376 50204
rect 183428 50192 183434 50244
rect 184842 50192 184848 50244
rect 184900 50232 184906 50244
rect 200666 50232 200672 50244
rect 184900 50204 200672 50232
rect 184900 50192 184906 50204
rect 200666 50192 200672 50204
rect 200724 50192 200730 50244
rect 201402 50192 201408 50244
rect 201460 50232 201466 50244
rect 214926 50232 214932 50244
rect 201460 50204 214932 50232
rect 201460 50192 201466 50204
rect 214926 50192 214932 50204
rect 214984 50192 214990 50244
rect 531866 50192 531872 50244
rect 531924 50232 531930 50244
rect 543001 50235 543059 50241
rect 543001 50232 543013 50235
rect 531924 50204 543013 50232
rect 531924 50192 531930 50204
rect 543001 50201 543013 50204
rect 543047 50201 543059 50235
rect 543001 50195 543059 50201
rect 88886 50164 88892 50176
rect 64846 50136 88892 50164
rect 88886 50124 88892 50136
rect 88944 50124 88950 50176
rect 88981 50167 89039 50173
rect 88981 50133 88993 50167
rect 89027 50164 89039 50167
rect 113266 50164 113272 50176
rect 89027 50136 113272 50164
rect 89027 50133 89039 50136
rect 88981 50127 89039 50133
rect 113266 50124 113272 50136
rect 113324 50124 113330 50176
rect 117222 50124 117228 50176
rect 117280 50164 117286 50176
rect 142798 50164 142804 50176
rect 117280 50136 142804 50164
rect 117280 50124 117286 50136
rect 142798 50124 142804 50136
rect 142856 50124 142862 50176
rect 150342 50124 150348 50176
rect 150400 50164 150406 50176
rect 171226 50164 171232 50176
rect 150400 50136 171232 50164
rect 150400 50124 150406 50136
rect 171226 50124 171232 50136
rect 171284 50124 171290 50176
rect 175182 50124 175188 50176
rect 175240 50164 175246 50176
rect 192570 50164 192576 50176
rect 175240 50136 192576 50164
rect 175240 50124 175246 50136
rect 192570 50124 192576 50136
rect 192628 50124 192634 50176
rect 195882 50124 195888 50176
rect 195940 50164 195946 50176
rect 210878 50164 210884 50176
rect 195940 50136 210884 50164
rect 195940 50124 195946 50136
rect 210878 50124 210884 50136
rect 210936 50124 210942 50176
rect 533890 50124 533896 50176
rect 533948 50164 533954 50176
rect 545758 50164 545764 50176
rect 533948 50136 545764 50164
rect 533948 50124 533954 50136
rect 545758 50124 545764 50136
rect 545816 50124 545822 50176
rect 35802 50056 35808 50108
rect 35860 50096 35866 50108
rect 72694 50096 72700 50108
rect 35860 50068 72700 50096
rect 35860 50056 35866 50068
rect 72694 50056 72700 50068
rect 72752 50056 72758 50108
rect 76742 50096 76748 50108
rect 74506 50068 76748 50096
rect 39942 49988 39948 50040
rect 40000 50028 40006 50040
rect 74506 50028 74534 50068
rect 76742 50056 76748 50068
rect 76800 50056 76806 50108
rect 78582 50056 78588 50108
rect 78640 50096 78646 50108
rect 81897 50099 81955 50105
rect 81897 50096 81909 50099
rect 78640 50068 81909 50096
rect 78640 50056 78646 50068
rect 81897 50065 81909 50068
rect 81943 50065 81955 50099
rect 81897 50059 81955 50065
rect 85482 50056 85488 50108
rect 85540 50096 85546 50108
rect 115382 50096 115388 50108
rect 85540 50068 115388 50096
rect 85540 50056 85546 50068
rect 115382 50056 115388 50068
rect 115440 50056 115446 50108
rect 118602 50056 118608 50108
rect 118660 50096 118666 50108
rect 143810 50096 143816 50108
rect 118660 50068 143816 50096
rect 118660 50056 118666 50068
rect 143810 50056 143816 50068
rect 143868 50056 143874 50108
rect 147582 50056 147588 50108
rect 147640 50096 147646 50108
rect 169202 50096 169208 50108
rect 147640 50068 169208 50096
rect 147640 50056 147646 50068
rect 169202 50056 169208 50068
rect 169260 50056 169266 50108
rect 176562 50056 176568 50108
rect 176620 50096 176626 50108
rect 193582 50096 193588 50108
rect 176620 50068 193588 50096
rect 176620 50056 176626 50068
rect 193582 50056 193588 50068
rect 193640 50056 193646 50108
rect 40000 50000 74534 50028
rect 40000 49988 40006 50000
rect 83458 49988 83464 50040
rect 83516 50028 83522 50040
rect 88981 50031 89039 50037
rect 88981 50028 88993 50031
rect 83516 50000 88993 50028
rect 83516 49988 83522 50000
rect 88981 49997 88993 50000
rect 89027 49997 89039 50031
rect 88981 49991 89039 49997
rect 89073 50031 89131 50037
rect 89073 49997 89085 50031
rect 89119 50028 89131 50031
rect 116394 50028 116400 50040
rect 89119 50000 116400 50028
rect 89119 49997 89131 50000
rect 89073 49991 89131 49997
rect 116394 49988 116400 50000
rect 116452 49988 116458 50040
rect 123849 50031 123907 50037
rect 123849 50028 123861 50031
rect 122806 50000 123861 50028
rect 45462 49920 45468 49972
rect 45520 49960 45526 49972
rect 80790 49960 80796 49972
rect 45520 49932 80796 49960
rect 45520 49920 45526 49932
rect 80790 49920 80796 49932
rect 80848 49920 80854 49972
rect 82078 49920 82084 49972
rect 82136 49960 82142 49972
rect 110230 49960 110236 49972
rect 82136 49932 110236 49960
rect 82136 49920 82142 49932
rect 110230 49920 110236 49932
rect 110288 49920 110294 49972
rect 119890 49920 119896 49972
rect 119948 49960 119954 49972
rect 122806 49960 122834 50000
rect 123849 49997 123861 50000
rect 123895 49997 123907 50031
rect 125413 50031 125471 50037
rect 125413 50028 125425 50031
rect 123849 49991 123907 49997
rect 123956 50000 125425 50028
rect 119948 49932 122834 49960
rect 119948 49920 119954 49932
rect 43438 49852 43444 49904
rect 43496 49892 43502 49904
rect 69658 49892 69664 49904
rect 43496 49864 69664 49892
rect 43496 49852 43502 49864
rect 69658 49852 69664 49864
rect 69716 49852 69722 49904
rect 71130 49852 71136 49904
rect 71188 49892 71194 49904
rect 73706 49892 73712 49904
rect 71188 49864 73712 49892
rect 71188 49852 71194 49864
rect 73706 49852 73712 49864
rect 73764 49852 73770 49904
rect 75178 49852 75184 49904
rect 75236 49892 75242 49904
rect 104158 49892 104164 49904
rect 75236 49864 104164 49892
rect 75236 49852 75242 49864
rect 104158 49852 104164 49864
rect 104216 49852 104222 49904
rect 106918 49852 106924 49904
rect 106976 49892 106982 49904
rect 123956 49892 123984 50000
rect 125413 49997 125425 50000
rect 125459 49997 125471 50031
rect 125413 49991 125471 49997
rect 125502 49988 125508 50040
rect 125560 50028 125566 50040
rect 149882 50028 149888 50040
rect 125560 50000 149888 50028
rect 125560 49988 125566 50000
rect 149882 49988 149888 50000
rect 149940 49988 149946 50040
rect 154482 49988 154488 50040
rect 154540 50028 154546 50040
rect 175274 50028 175280 50040
rect 154540 50000 175280 50028
rect 154540 49988 154546 50000
rect 175274 49988 175280 50000
rect 175332 49988 175338 50040
rect 177942 49988 177948 50040
rect 178000 50028 178006 50040
rect 195606 50028 195612 50040
rect 178000 50000 195612 50028
rect 178000 49988 178006 50000
rect 195606 49988 195612 50000
rect 195664 49988 195670 50040
rect 263502 49988 263508 50040
rect 263560 50028 263566 50040
rect 268746 50028 268752 50040
rect 263560 50000 268752 50028
rect 263560 49988 263566 50000
rect 268746 49988 268752 50000
rect 268804 49988 268810 50040
rect 124033 49963 124091 49969
rect 124033 49929 124045 49963
rect 124079 49960 124091 49963
rect 144822 49960 144828 49972
rect 124079 49932 144828 49960
rect 124079 49929 124091 49932
rect 124033 49923 124091 49929
rect 144822 49920 144828 49932
rect 144880 49920 144886 49972
rect 151722 49920 151728 49972
rect 151780 49960 151786 49972
rect 172238 49960 172244 49972
rect 151780 49932 172244 49960
rect 151780 49920 151786 49932
rect 172238 49920 172244 49932
rect 172296 49920 172302 49972
rect 172333 49963 172391 49969
rect 172333 49929 172345 49963
rect 172379 49960 172391 49963
rect 172379 49932 173388 49960
rect 172379 49929 172391 49932
rect 172333 49923 172391 49929
rect 125134 49892 125140 49904
rect 106976 49864 123984 49892
rect 124048 49864 125140 49892
rect 106976 49852 106982 49864
rect 44818 49784 44824 49836
rect 44876 49824 44882 49836
rect 60458 49824 60464 49836
rect 44876 49796 60464 49824
rect 44876 49784 44882 49796
rect 60458 49784 60464 49796
rect 60516 49784 60522 49836
rect 64230 49784 64236 49836
rect 64288 49824 64294 49836
rect 64288 49796 84194 49824
rect 64288 49784 64294 49796
rect 46198 49716 46204 49768
rect 46256 49756 46262 49768
rect 47302 49756 47308 49768
rect 46256 49728 47308 49756
rect 46256 49716 46262 49728
rect 47302 49716 47308 49728
rect 47360 49716 47366 49768
rect 50338 49716 50344 49768
rect 50396 49756 50402 49768
rect 75730 49756 75736 49768
rect 50396 49728 75736 49756
rect 50396 49716 50402 49728
rect 75730 49716 75736 49728
rect 75788 49716 75794 49768
rect 76558 49716 76564 49768
rect 76616 49756 76622 49768
rect 82814 49756 82820 49768
rect 76616 49728 82820 49756
rect 76616 49716 76622 49728
rect 82814 49716 82820 49728
rect 82872 49716 82878 49768
rect 84166 49756 84194 49796
rect 86862 49784 86868 49836
rect 86920 49824 86926 49836
rect 89073 49827 89131 49833
rect 89073 49824 89085 49827
rect 86920 49796 89085 49824
rect 86920 49784 86926 49796
rect 89073 49793 89085 49796
rect 89119 49793 89131 49827
rect 89073 49787 89131 49793
rect 95878 49784 95884 49836
rect 95936 49824 95942 49836
rect 122466 49824 122472 49836
rect 95936 49796 122472 49824
rect 95936 49784 95942 49796
rect 122466 49784 122472 49796
rect 122524 49784 122530 49836
rect 92014 49756 92020 49768
rect 84166 49728 92020 49756
rect 92014 49716 92020 49728
rect 92072 49716 92078 49768
rect 93118 49716 93124 49768
rect 93176 49756 93182 49768
rect 98086 49756 98092 49768
rect 93176 49728 98092 49756
rect 93176 49716 93182 49728
rect 98086 49716 98092 49728
rect 98144 49716 98150 49768
rect 98638 49716 98644 49768
rect 98696 49756 98702 49768
rect 124048 49756 124076 49864
rect 125134 49852 125140 49864
rect 125192 49852 125198 49904
rect 140774 49892 140780 49904
rect 134536 49864 140780 49892
rect 124122 49784 124128 49836
rect 124180 49824 124186 49836
rect 134337 49827 134395 49833
rect 134337 49824 134349 49827
rect 124180 49796 134349 49824
rect 124180 49784 124186 49796
rect 134337 49793 134349 49796
rect 134383 49793 134395 49827
rect 134337 49787 134395 49793
rect 98696 49728 124076 49756
rect 98696 49716 98702 49728
rect 124858 49716 124864 49768
rect 124916 49756 124922 49768
rect 134536 49756 134564 49864
rect 140774 49852 140780 49864
rect 140832 49852 140838 49904
rect 146202 49852 146208 49904
rect 146260 49892 146266 49904
rect 153013 49895 153071 49901
rect 153013 49892 153025 49895
rect 146260 49864 153025 49892
rect 146260 49852 146266 49864
rect 153013 49861 153025 49864
rect 153059 49861 153071 49895
rect 153013 49855 153071 49861
rect 153102 49852 153108 49904
rect 153160 49892 153166 49904
rect 173250 49892 173256 49904
rect 153160 49864 173256 49892
rect 153160 49852 153166 49864
rect 173250 49852 173256 49864
rect 173308 49852 173314 49904
rect 173360 49892 173388 49932
rect 173802 49920 173808 49972
rect 173860 49960 173866 49972
rect 191558 49960 191564 49972
rect 173860 49932 191564 49960
rect 173860 49920 173866 49932
rect 191558 49920 191564 49932
rect 191616 49920 191622 49972
rect 193122 49920 193128 49972
rect 193180 49960 193186 49972
rect 207750 49960 207756 49972
rect 193180 49932 207756 49960
rect 193180 49920 193186 49932
rect 207750 49920 207756 49932
rect 207808 49920 207814 49972
rect 270402 49920 270408 49972
rect 270460 49960 270466 49972
rect 274818 49960 274824 49972
rect 270460 49932 274824 49960
rect 270460 49920 270466 49932
rect 274818 49920 274824 49932
rect 274876 49920 274882 49972
rect 177298 49892 177304 49904
rect 173360 49864 177304 49892
rect 177298 49852 177304 49864
rect 177356 49852 177362 49904
rect 182082 49852 182088 49904
rect 182140 49892 182146 49904
rect 198366 49892 198372 49904
rect 182140 49864 198372 49892
rect 182140 49852 182146 49864
rect 198366 49852 198372 49864
rect 198424 49852 198430 49904
rect 260650 49852 260656 49904
rect 260708 49892 260714 49904
rect 266722 49892 266728 49904
rect 260708 49864 266728 49892
rect 260708 49852 260714 49864
rect 266722 49852 266728 49864
rect 266780 49852 266786 49904
rect 269022 49852 269028 49904
rect 269080 49892 269086 49904
rect 273806 49892 273812 49904
rect 269080 49864 273812 49892
rect 269080 49852 269086 49864
rect 273806 49852 273812 49864
rect 273864 49852 273870 49904
rect 280062 49852 280068 49904
rect 280120 49892 280126 49904
rect 283006 49892 283012 49904
rect 280120 49864 283012 49892
rect 280120 49852 280126 49864
rect 283006 49852 283012 49864
rect 283064 49852 283070 49904
rect 313458 49852 313464 49904
rect 313516 49892 313522 49904
rect 314470 49892 314476 49904
rect 313516 49864 314476 49892
rect 313516 49852 313522 49864
rect 314470 49852 314476 49864
rect 314528 49852 314534 49904
rect 513558 49852 513564 49904
rect 513616 49892 513622 49904
rect 519538 49892 519544 49904
rect 513616 49864 519544 49892
rect 513616 49852 513622 49864
rect 519538 49852 519544 49864
rect 519596 49852 519602 49904
rect 540974 49852 540980 49904
rect 541032 49892 541038 49904
rect 548610 49892 548616 49904
rect 541032 49864 548616 49892
rect 541032 49852 541038 49864
rect 548610 49852 548616 49864
rect 548668 49852 548674 49904
rect 134613 49827 134671 49833
rect 134613 49793 134625 49827
rect 134659 49824 134671 49827
rect 148870 49824 148876 49836
rect 134659 49796 148876 49824
rect 134659 49793 134671 49796
rect 134613 49787 134671 49793
rect 148870 49784 148876 49796
rect 148928 49784 148934 49836
rect 155862 49784 155868 49836
rect 155920 49824 155926 49836
rect 176286 49824 176292 49836
rect 155920 49796 176292 49824
rect 155920 49784 155926 49796
rect 176286 49784 176292 49796
rect 176344 49784 176350 49836
rect 249702 49784 249708 49836
rect 249760 49824 249766 49836
rect 256510 49824 256516 49836
rect 249760 49796 256516 49824
rect 249760 49784 249766 49796
rect 256510 49784 256516 49796
rect 256568 49784 256574 49836
rect 259362 49784 259368 49836
rect 259420 49824 259426 49836
rect 264698 49824 264704 49836
rect 259420 49796 264704 49824
rect 259420 49784 259426 49796
rect 264698 49784 264704 49796
rect 264756 49784 264762 49836
rect 271782 49784 271788 49836
rect 271840 49824 271846 49836
rect 275830 49824 275836 49836
rect 271840 49796 275836 49824
rect 271840 49784 271846 49796
rect 275830 49784 275836 49796
rect 275888 49784 275894 49836
rect 281442 49784 281448 49836
rect 281500 49824 281506 49836
rect 284018 49824 284024 49836
rect 281500 49796 284024 49824
rect 281500 49784 281506 49796
rect 284018 49784 284024 49796
rect 284076 49784 284082 49836
rect 288342 49784 288348 49836
rect 288400 49824 288406 49836
rect 290090 49824 290096 49836
rect 288400 49796 290096 49824
rect 288400 49784 288406 49796
rect 290090 49784 290096 49796
rect 290148 49784 290154 49836
rect 317506 49784 317512 49836
rect 317564 49824 317570 49836
rect 318702 49824 318708 49836
rect 317564 49796 318708 49824
rect 317564 49784 317570 49796
rect 318702 49784 318708 49796
rect 318760 49784 318766 49836
rect 319530 49784 319536 49836
rect 319588 49824 319594 49836
rect 320818 49824 320824 49836
rect 319588 49796 320824 49824
rect 319588 49784 319594 49796
rect 320818 49784 320824 49796
rect 320876 49784 320882 49836
rect 336826 49784 336832 49836
rect 336884 49824 336890 49836
rect 338850 49824 338856 49836
rect 336884 49796 338856 49824
rect 336884 49784 336890 49796
rect 338850 49784 338856 49796
rect 338908 49784 338914 49836
rect 434346 49784 434352 49836
rect 434404 49824 434410 49836
rect 435358 49824 435364 49836
rect 434404 49796 435364 49824
rect 434404 49784 434410 49796
rect 435358 49784 435364 49796
rect 435416 49784 435422 49836
rect 451642 49784 451648 49836
rect 451700 49824 451706 49836
rect 454678 49824 454684 49836
rect 451700 49796 454684 49824
rect 451700 49784 451706 49796
rect 454678 49784 454684 49796
rect 454736 49784 454742 49836
rect 124916 49728 134564 49756
rect 124916 49716 124922 49728
rect 137278 49716 137284 49768
rect 137336 49756 137342 49768
rect 138750 49756 138756 49768
rect 137336 49728 138756 49756
rect 137336 49716 137342 49728
rect 138750 49716 138756 49728
rect 138808 49716 138814 49768
rect 157242 49716 157248 49768
rect 157300 49756 157306 49768
rect 172333 49759 172391 49765
rect 172333 49756 172345 49759
rect 157300 49728 172345 49756
rect 157300 49716 157306 49728
rect 172333 49725 172345 49728
rect 172379 49725 172391 49759
rect 172333 49719 172391 49725
rect 172422 49716 172428 49768
rect 172480 49756 172486 49768
rect 180521 49759 180579 49765
rect 180521 49756 180533 49759
rect 172480 49728 180533 49756
rect 172480 49716 172486 49728
rect 180521 49725 180533 49728
rect 180567 49725 180579 49759
rect 180521 49719 180579 49725
rect 251082 49716 251088 49768
rect 251140 49756 251146 49768
rect 257522 49756 257528 49768
rect 251140 49728 257528 49756
rect 251140 49716 251146 49728
rect 257522 49716 257528 49728
rect 257580 49716 257586 49768
rect 260742 49716 260748 49768
rect 260800 49756 260806 49768
rect 265710 49756 265716 49768
rect 260800 49728 265716 49756
rect 260800 49716 260806 49728
rect 265710 49716 265716 49728
rect 265768 49716 265774 49768
rect 268930 49716 268936 49768
rect 268988 49756 268994 49768
rect 272794 49756 272800 49768
rect 268988 49728 272800 49756
rect 268988 49716 268994 49728
rect 272794 49716 272800 49728
rect 272852 49716 272858 49768
rect 273898 49716 273904 49768
rect 273956 49756 273962 49768
rect 276842 49756 276848 49768
rect 273956 49728 276848 49756
rect 273956 49716 273962 49728
rect 276842 49716 276848 49728
rect 276900 49716 276906 49768
rect 278682 49716 278688 49768
rect 278740 49756 278746 49768
rect 281994 49756 282000 49768
rect 278740 49728 282000 49756
rect 278740 49716 278746 49728
rect 281994 49716 282000 49728
rect 282052 49716 282058 49768
rect 282822 49716 282828 49768
rect 282880 49756 282886 49768
rect 285030 49756 285036 49768
rect 282880 49728 285036 49756
rect 282880 49716 282886 49728
rect 285030 49716 285036 49728
rect 285088 49716 285094 49768
rect 289722 49716 289728 49768
rect 289780 49756 289786 49768
rect 291102 49756 291108 49768
rect 289780 49728 291108 49756
rect 289780 49716 289786 49728
rect 291102 49716 291108 49728
rect 291160 49716 291166 49768
rect 312446 49716 312452 49768
rect 312504 49756 312510 49768
rect 313458 49756 313464 49768
rect 312504 49728 313464 49756
rect 312504 49716 312510 49728
rect 313458 49716 313464 49728
rect 313516 49716 313522 49768
rect 316494 49716 316500 49768
rect 316552 49756 316558 49768
rect 317598 49756 317604 49768
rect 316552 49728 317604 49756
rect 316552 49716 316558 49728
rect 317598 49716 317604 49728
rect 317656 49716 317662 49768
rect 320542 49716 320548 49768
rect 320600 49756 320606 49768
rect 321462 49756 321468 49768
rect 320600 49728 321468 49756
rect 320600 49716 320606 49728
rect 321462 49716 321468 49728
rect 321520 49716 321526 49768
rect 321554 49716 321560 49768
rect 321612 49756 321618 49768
rect 322750 49756 322756 49768
rect 321612 49728 322756 49756
rect 321612 49716 321618 49728
rect 322750 49716 322756 49728
rect 322808 49716 322814 49768
rect 324590 49716 324596 49768
rect 324648 49756 324654 49768
rect 325510 49756 325516 49768
rect 324648 49728 325516 49756
rect 324648 49716 324654 49728
rect 325510 49716 325516 49728
rect 325568 49716 325574 49768
rect 328638 49716 328644 49768
rect 328696 49756 328702 49768
rect 329742 49756 329748 49768
rect 328696 49728 329748 49756
rect 328696 49716 328702 49728
rect 329742 49716 329748 49728
rect 329800 49716 329806 49768
rect 331766 49716 331772 49768
rect 331824 49756 331830 49768
rect 332502 49756 332508 49768
rect 331824 49728 332508 49756
rect 331824 49716 331830 49728
rect 332502 49716 332508 49728
rect 332560 49716 332566 49768
rect 333790 49716 333796 49768
rect 333848 49756 333854 49768
rect 334618 49756 334624 49768
rect 333848 49728 334624 49756
rect 333848 49716 333854 49728
rect 334618 49716 334624 49728
rect 334676 49716 334682 49768
rect 335814 49716 335820 49768
rect 335872 49756 335878 49768
rect 336642 49756 336648 49768
rect 335872 49728 336648 49756
rect 335872 49716 335878 49728
rect 336642 49716 336648 49728
rect 336700 49716 336706 49768
rect 337838 49716 337844 49768
rect 337896 49756 337902 49768
rect 338758 49756 338764 49768
rect 337896 49728 338764 49756
rect 337896 49716 337902 49728
rect 338758 49716 338764 49728
rect 338816 49716 338822 49768
rect 339862 49716 339868 49768
rect 339920 49756 339926 49768
rect 340782 49756 340788 49768
rect 339920 49728 340788 49756
rect 339920 49716 339926 49728
rect 340782 49716 340788 49728
rect 340840 49716 340846 49768
rect 340874 49716 340880 49768
rect 340932 49756 340938 49768
rect 342162 49756 342168 49768
rect 340932 49728 342168 49756
rect 340932 49716 340938 49728
rect 342162 49716 342168 49728
rect 342220 49716 342226 49768
rect 347958 49716 347964 49768
rect 348016 49756 348022 49768
rect 348970 49756 348976 49768
rect 348016 49728 348976 49756
rect 348016 49716 348022 49728
rect 348970 49716 348976 49728
rect 349028 49716 349034 49768
rect 350994 49716 351000 49768
rect 351052 49756 351058 49768
rect 351822 49756 351828 49768
rect 351052 49728 351828 49756
rect 351052 49716 351058 49728
rect 351822 49716 351828 49728
rect 351880 49716 351886 49768
rect 352006 49716 352012 49768
rect 352064 49756 352070 49768
rect 353110 49756 353116 49768
rect 352064 49728 353116 49756
rect 352064 49716 352070 49728
rect 353110 49716 353116 49728
rect 353168 49716 353174 49768
rect 355134 49716 355140 49768
rect 355192 49756 355198 49768
rect 355962 49756 355968 49768
rect 355192 49728 355968 49756
rect 355192 49716 355198 49728
rect 355962 49716 355968 49728
rect 356020 49716 356026 49768
rect 356146 49716 356152 49768
rect 356204 49756 356210 49768
rect 357342 49756 357348 49768
rect 356204 49728 357348 49756
rect 356204 49716 356210 49728
rect 357342 49716 357348 49728
rect 357400 49716 357406 49768
rect 359182 49716 359188 49768
rect 359240 49756 359246 49768
rect 360102 49756 360108 49768
rect 359240 49728 360108 49756
rect 359240 49716 359246 49728
rect 360102 49716 360108 49728
rect 360160 49716 360166 49768
rect 360194 49716 360200 49768
rect 360252 49756 360258 49768
rect 361482 49756 361488 49768
rect 360252 49728 361488 49756
rect 360252 49716 360258 49728
rect 361482 49716 361488 49728
rect 361540 49716 361546 49768
rect 363230 49716 363236 49768
rect 363288 49756 363294 49768
rect 364150 49756 364156 49768
rect 363288 49728 364156 49756
rect 363288 49716 363294 49728
rect 364150 49716 364156 49728
rect 364208 49716 364214 49768
rect 367278 49716 367284 49768
rect 367336 49756 367342 49768
rect 368290 49756 368296 49768
rect 367336 49728 368296 49756
rect 367336 49716 367342 49728
rect 368290 49716 368296 49728
rect 368348 49716 368354 49768
rect 370314 49716 370320 49768
rect 370372 49756 370378 49768
rect 371142 49756 371148 49768
rect 370372 49728 371148 49756
rect 370372 49716 370378 49728
rect 371142 49716 371148 49728
rect 371200 49716 371206 49768
rect 371326 49716 371332 49768
rect 371384 49756 371390 49768
rect 372522 49756 372528 49768
rect 371384 49728 372528 49756
rect 371384 49716 371390 49728
rect 372522 49716 372528 49728
rect 372580 49716 372586 49768
rect 374362 49716 374368 49768
rect 374420 49756 374426 49768
rect 375282 49756 375288 49768
rect 374420 49728 375288 49756
rect 374420 49716 374426 49728
rect 375282 49716 375288 49728
rect 375340 49716 375346 49768
rect 375374 49716 375380 49768
rect 375432 49756 375438 49768
rect 376570 49756 376576 49768
rect 375432 49728 376576 49756
rect 375432 49716 375438 49728
rect 376570 49716 376576 49728
rect 376628 49716 376634 49768
rect 378502 49716 378508 49768
rect 378560 49756 378566 49768
rect 379422 49756 379428 49768
rect 378560 49728 379428 49756
rect 378560 49716 378566 49728
rect 379422 49716 379428 49728
rect 379480 49716 379486 49768
rect 379514 49716 379520 49768
rect 379572 49756 379578 49768
rect 380710 49756 380716 49768
rect 379572 49728 380716 49756
rect 379572 49716 379578 49728
rect 380710 49716 380716 49728
rect 380768 49716 380774 49768
rect 382550 49716 382556 49768
rect 382608 49756 382614 49768
rect 383470 49756 383476 49768
rect 382608 49728 383476 49756
rect 382608 49716 382614 49728
rect 383470 49716 383476 49728
rect 383528 49716 383534 49768
rect 386598 49716 386604 49768
rect 386656 49756 386662 49768
rect 387702 49756 387708 49768
rect 386656 49728 387708 49756
rect 386656 49716 386662 49728
rect 387702 49716 387708 49728
rect 387760 49716 387766 49768
rect 389634 49716 389640 49768
rect 389692 49756 389698 49768
rect 390462 49756 390468 49768
rect 389692 49728 390468 49756
rect 389692 49716 389698 49728
rect 390462 49716 390468 49728
rect 390520 49716 390526 49768
rect 390646 49716 390652 49768
rect 390704 49756 390710 49768
rect 391750 49756 391756 49768
rect 390704 49728 391756 49756
rect 390704 49716 390710 49728
rect 391750 49716 391756 49728
rect 391808 49716 391814 49768
rect 393682 49716 393688 49768
rect 393740 49756 393746 49768
rect 394602 49756 394608 49768
rect 393740 49728 394608 49756
rect 393740 49716 393746 49728
rect 394602 49716 394608 49728
rect 394660 49716 394666 49768
rect 394694 49716 394700 49768
rect 394752 49756 394758 49768
rect 395890 49756 395896 49768
rect 394752 49728 395896 49756
rect 394752 49716 394758 49728
rect 395890 49716 395896 49728
rect 395948 49716 395954 49768
rect 397730 49716 397736 49768
rect 397788 49756 397794 49768
rect 398650 49756 398656 49768
rect 397788 49728 398656 49756
rect 397788 49716 397794 49728
rect 398650 49716 398656 49728
rect 398708 49716 398714 49768
rect 400766 49716 400772 49768
rect 400824 49756 400830 49768
rect 401502 49756 401508 49768
rect 400824 49728 401508 49756
rect 400824 49716 400830 49728
rect 401502 49716 401508 49728
rect 401560 49716 401566 49768
rect 401870 49716 401876 49768
rect 401928 49756 401934 49768
rect 402882 49756 402888 49768
rect 401928 49728 402888 49756
rect 401928 49716 401934 49728
rect 402882 49716 402888 49728
rect 402940 49716 402946 49768
rect 405918 49716 405924 49768
rect 405976 49756 405982 49768
rect 406930 49756 406936 49768
rect 405976 49728 406936 49756
rect 405976 49716 405982 49728
rect 406930 49716 406936 49728
rect 406988 49716 406994 49768
rect 408954 49716 408960 49768
rect 409012 49756 409018 49768
rect 409782 49756 409788 49768
rect 409012 49728 409788 49756
rect 409012 49716 409018 49728
rect 409782 49716 409788 49728
rect 409840 49716 409846 49768
rect 409966 49716 409972 49768
rect 410024 49756 410030 49768
rect 411070 49756 411076 49768
rect 410024 49728 411076 49756
rect 410024 49716 410030 49728
rect 411070 49716 411076 49728
rect 411128 49716 411134 49768
rect 413002 49716 413008 49768
rect 413060 49756 413066 49768
rect 413922 49756 413928 49768
rect 413060 49728 413928 49756
rect 413060 49716 413066 49728
rect 413922 49716 413928 49728
rect 413980 49716 413986 49768
rect 414014 49716 414020 49768
rect 414072 49756 414078 49768
rect 415302 49756 415308 49768
rect 414072 49728 415308 49756
rect 414072 49716 414078 49728
rect 415302 49716 415308 49728
rect 415360 49716 415366 49768
rect 417050 49716 417056 49768
rect 417108 49756 417114 49768
rect 418062 49756 418068 49768
rect 417108 49728 418068 49756
rect 417108 49716 417114 49728
rect 418062 49716 418068 49728
rect 418120 49716 418126 49768
rect 420086 49716 420092 49768
rect 420144 49756 420150 49768
rect 420822 49756 420828 49768
rect 420144 49728 420828 49756
rect 420144 49716 420150 49728
rect 420822 49716 420828 49728
rect 420880 49716 420886 49768
rect 421098 49716 421104 49768
rect 421156 49756 421162 49768
rect 422202 49756 422208 49768
rect 421156 49728 422208 49756
rect 421156 49716 421162 49728
rect 422202 49716 422208 49728
rect 422260 49716 422266 49768
rect 424134 49716 424140 49768
rect 424192 49756 424198 49768
rect 424962 49756 424968 49768
rect 424192 49728 424968 49756
rect 424192 49716 424198 49728
rect 424962 49716 424968 49728
rect 425020 49716 425026 49768
rect 425238 49716 425244 49768
rect 425296 49756 425302 49768
rect 426250 49756 426256 49768
rect 425296 49728 426256 49756
rect 425296 49716 425302 49728
rect 426250 49716 426256 49728
rect 426308 49716 426314 49768
rect 428274 49716 428280 49768
rect 428332 49756 428338 49768
rect 429102 49756 429108 49768
rect 428332 49728 429108 49756
rect 428332 49716 428338 49728
rect 429102 49716 429108 49728
rect 429160 49716 429166 49768
rect 429286 49716 429292 49768
rect 429344 49756 429350 49768
rect 430482 49756 430488 49768
rect 429344 49728 430488 49756
rect 429344 49716 429350 49728
rect 430482 49716 430488 49728
rect 430540 49716 430546 49768
rect 432322 49716 432328 49768
rect 432380 49756 432386 49768
rect 433242 49756 433248 49768
rect 432380 49728 433248 49756
rect 432380 49716 432386 49728
rect 433242 49716 433248 49728
rect 433300 49716 433306 49768
rect 433334 49716 433340 49768
rect 433392 49756 433398 49768
rect 434622 49756 434628 49768
rect 433392 49728 434628 49756
rect 433392 49716 433398 49728
rect 434622 49716 434628 49728
rect 434680 49716 434686 49768
rect 436370 49716 436376 49768
rect 436428 49756 436434 49768
rect 437382 49756 437388 49768
rect 436428 49728 437388 49756
rect 436428 49716 436434 49728
rect 437382 49716 437388 49728
rect 437440 49716 437446 49768
rect 439406 49716 439412 49768
rect 439464 49756 439470 49768
rect 440142 49756 440148 49768
rect 439464 49728 440148 49756
rect 439464 49716 439470 49728
rect 440142 49716 440148 49728
rect 440200 49716 440206 49768
rect 443454 49716 443460 49768
rect 443512 49756 443518 49768
rect 444282 49756 444288 49768
rect 443512 49728 444288 49756
rect 443512 49716 443518 49728
rect 444282 49716 444288 49728
rect 444340 49716 444346 49768
rect 444466 49716 444472 49768
rect 444524 49756 444530 49768
rect 445662 49756 445668 49768
rect 444524 49728 445668 49756
rect 444524 49716 444530 49728
rect 445662 49716 445668 49728
rect 445720 49716 445726 49768
rect 447502 49716 447508 49768
rect 447560 49756 447566 49768
rect 448422 49756 448428 49768
rect 447560 49728 448428 49756
rect 447560 49716 447566 49728
rect 448422 49716 448428 49728
rect 448480 49716 448486 49768
rect 448514 49716 448520 49768
rect 448572 49756 448578 49768
rect 449802 49756 449808 49768
rect 448572 49728 449808 49756
rect 448572 49716 448578 49728
rect 449802 49716 449808 49728
rect 449860 49716 449866 49768
rect 452654 49716 452660 49768
rect 452712 49756 452718 49768
rect 453850 49756 453856 49768
rect 452712 49728 453856 49756
rect 452712 49716 452718 49728
rect 453850 49716 453856 49728
rect 453908 49716 453914 49768
rect 455690 49716 455696 49768
rect 455748 49756 455754 49768
rect 457438 49756 457444 49768
rect 455748 49728 457444 49756
rect 455748 49716 455754 49728
rect 457438 49716 457444 49728
rect 457496 49716 457502 49768
rect 459738 49716 459744 49768
rect 459796 49756 459802 49768
rect 460750 49756 460756 49768
rect 459796 49728 460756 49756
rect 459796 49716 459802 49728
rect 460750 49716 460756 49728
rect 460808 49716 460814 49768
rect 462774 49716 462780 49768
rect 462832 49756 462838 49768
rect 463602 49756 463608 49768
rect 462832 49728 463608 49756
rect 462832 49716 462838 49728
rect 463602 49716 463608 49728
rect 463660 49716 463666 49768
rect 463786 49716 463792 49768
rect 463844 49756 463850 49768
rect 464982 49756 464988 49768
rect 463844 49728 464988 49756
rect 463844 49716 463850 49728
rect 464982 49716 464988 49728
rect 465040 49716 465046 49768
rect 466822 49716 466828 49768
rect 466880 49756 466886 49768
rect 467742 49756 467748 49768
rect 466880 49728 467748 49756
rect 466880 49716 466886 49728
rect 467742 49716 467748 49728
rect 467800 49716 467806 49768
rect 467834 49716 467840 49768
rect 467892 49756 467898 49768
rect 469030 49756 469036 49768
rect 467892 49728 469036 49756
rect 467892 49716 467898 49728
rect 469030 49716 469036 49728
rect 469088 49716 469094 49768
rect 470870 49716 470876 49768
rect 470928 49756 470934 49768
rect 471790 49756 471796 49768
rect 470928 49728 471796 49756
rect 470928 49716 470934 49728
rect 471790 49716 471796 49728
rect 471848 49716 471854 49768
rect 475010 49716 475016 49768
rect 475068 49756 475074 49768
rect 475930 49756 475936 49768
rect 475068 49728 475936 49756
rect 475068 49716 475074 49728
rect 475930 49716 475936 49728
rect 475988 49716 475994 49768
rect 478046 49716 478052 49768
rect 478104 49756 478110 49768
rect 478782 49756 478788 49768
rect 478104 49728 478788 49756
rect 478104 49716 478110 49728
rect 478782 49716 478788 49728
rect 478840 49716 478846 49768
rect 479058 49716 479064 49768
rect 479116 49756 479122 49768
rect 480162 49756 480168 49768
rect 479116 49728 480168 49756
rect 479116 49716 479122 49728
rect 480162 49716 480168 49728
rect 480220 49716 480226 49768
rect 482094 49716 482100 49768
rect 482152 49756 482158 49768
rect 482922 49756 482928 49768
rect 482152 49728 482928 49756
rect 482152 49716 482158 49728
rect 482922 49716 482928 49728
rect 482980 49716 482986 49768
rect 483106 49716 483112 49768
rect 483164 49756 483170 49768
rect 484210 49756 484216 49768
rect 483164 49728 484216 49756
rect 483164 49716 483170 49728
rect 484210 49716 484216 49728
rect 484268 49716 484274 49768
rect 486142 49716 486148 49768
rect 486200 49756 486206 49768
rect 487062 49756 487068 49768
rect 486200 49728 487068 49756
rect 486200 49716 486206 49728
rect 487062 49716 487068 49728
rect 487120 49716 487126 49768
rect 487154 49716 487160 49768
rect 487212 49756 487218 49768
rect 488442 49756 488448 49768
rect 487212 49728 488448 49756
rect 487212 49716 487218 49728
rect 488442 49716 488448 49728
rect 488500 49716 488506 49768
rect 490190 49716 490196 49768
rect 490248 49756 490254 49768
rect 491110 49756 491116 49768
rect 490248 49728 491116 49756
rect 490248 49716 490254 49728
rect 491110 49716 491116 49728
rect 491168 49716 491174 49768
rect 497366 49716 497372 49768
rect 497424 49756 497430 49768
rect 498102 49756 498108 49768
rect 497424 49728 498108 49756
rect 497424 49716 497430 49728
rect 498102 49716 498108 49728
rect 498160 49716 498166 49768
rect 501414 49716 501420 49768
rect 501472 49756 501478 49768
rect 502242 49756 502248 49768
rect 501472 49728 502248 49756
rect 501472 49716 501478 49728
rect 502242 49716 502248 49728
rect 502300 49716 502306 49768
rect 502426 49716 502432 49768
rect 502484 49756 502490 49768
rect 503622 49756 503628 49768
rect 502484 49728 503628 49756
rect 502484 49716 502490 49728
rect 503622 49716 503628 49728
rect 503680 49716 503686 49768
rect 505462 49716 505468 49768
rect 505520 49756 505526 49768
rect 506382 49756 506388 49768
rect 505520 49728 506388 49756
rect 505520 49716 505526 49728
rect 506382 49716 506388 49728
rect 506440 49716 506446 49768
rect 517606 49716 517612 49768
rect 517664 49756 517670 49768
rect 518710 49756 518716 49768
rect 517664 49728 518716 49756
rect 517664 49716 517670 49728
rect 518710 49716 518716 49728
rect 518768 49716 518774 49768
rect 520734 49716 520740 49768
rect 520792 49756 520798 49768
rect 521562 49756 521568 49768
rect 520792 49728 521568 49756
rect 520792 49716 520798 49728
rect 521562 49716 521568 49728
rect 521620 49716 521626 49768
rect 521746 49716 521752 49768
rect 521804 49756 521810 49768
rect 522942 49756 522948 49768
rect 521804 49728 522948 49756
rect 521804 49716 521810 49728
rect 522942 49716 522948 49728
rect 523000 49716 523006 49768
rect 524782 49716 524788 49768
rect 524840 49756 524846 49768
rect 525702 49756 525708 49768
rect 524840 49728 525708 49756
rect 524840 49716 524846 49728
rect 525702 49716 525708 49728
rect 525760 49716 525766 49768
rect 532878 49716 532884 49768
rect 532936 49756 532942 49768
rect 533982 49756 533988 49768
rect 532936 49728 533988 49756
rect 532936 49716 532942 49728
rect 533982 49716 533988 49728
rect 534040 49716 534046 49768
rect 535914 49716 535920 49768
rect 535972 49756 535978 49768
rect 536742 49756 536748 49768
rect 535972 49728 536748 49756
rect 535972 49716 535978 49728
rect 536742 49716 536748 49728
rect 536800 49716 536806 49768
rect 536926 49716 536932 49768
rect 536984 49756 536990 49768
rect 538122 49756 538128 49768
rect 536984 49728 538128 49756
rect 536984 49716 536990 49728
rect 538122 49716 538128 49728
rect 538180 49716 538186 49768
rect 539962 49716 539968 49768
rect 540020 49756 540026 49768
rect 547138 49756 547144 49768
rect 540020 49728 547144 49756
rect 540020 49716 540026 49728
rect 547138 49716 547144 49728
rect 547196 49716 547202 49768
rect 66162 49580 66168 49632
rect 66220 49620 66226 49632
rect 99098 49620 99104 49632
rect 66220 49592 99104 49620
rect 66220 49580 66226 49592
rect 99098 49580 99104 49592
rect 99156 49580 99162 49632
rect 70210 49512 70216 49564
rect 70268 49552 70274 49564
rect 102134 49552 102140 49564
rect 70268 49524 102140 49552
rect 70268 49512 70274 49524
rect 102134 49512 102140 49524
rect 102192 49512 102198 49564
rect 41322 49444 41328 49496
rect 41380 49484 41386 49496
rect 77202 49484 77208 49496
rect 41380 49456 77208 49484
rect 41380 49444 41386 49456
rect 77202 49444 77208 49456
rect 77260 49444 77266 49496
rect 84102 49444 84108 49496
rect 84160 49484 84166 49496
rect 114278 49484 114284 49496
rect 84160 49456 114284 49484
rect 84160 49444 84166 49456
rect 114278 49444 114284 49456
rect 114336 49444 114342 49496
rect 34422 49376 34428 49428
rect 34480 49416 34486 49428
rect 71682 49416 71688 49428
rect 34480 49388 71688 49416
rect 34480 49376 34486 49388
rect 71682 49376 71688 49388
rect 71740 49376 71746 49428
rect 73062 49376 73068 49428
rect 73120 49416 73126 49428
rect 105170 49416 105176 49428
rect 73120 49388 105176 49416
rect 73120 49376 73126 49388
rect 105170 49376 105176 49388
rect 105228 49376 105234 49428
rect 7558 49308 7564 49360
rect 7616 49348 7622 49360
rect 44266 49348 44272 49360
rect 7616 49320 44272 49348
rect 7616 49308 7622 49320
rect 44266 49308 44272 49320
rect 44324 49308 44330 49360
rect 52362 49308 52368 49360
rect 52420 49348 52426 49360
rect 86494 49348 86500 49360
rect 52420 49320 86500 49348
rect 52420 49308 52426 49320
rect 86494 49308 86500 49320
rect 86552 49308 86558 49360
rect 102042 49308 102048 49360
rect 102100 49348 102106 49360
rect 129550 49348 129556 49360
rect 102100 49320 129556 49348
rect 102100 49308 102106 49320
rect 129550 49308 129556 49320
rect 129608 49308 129614 49360
rect 298094 49308 298100 49360
rect 298152 49348 298158 49360
rect 298830 49348 298836 49360
rect 298152 49320 298836 49348
rect 298152 49308 298158 49320
rect 298830 49308 298836 49320
rect 298888 49308 298894 49360
rect 37182 49240 37188 49292
rect 37240 49280 37246 49292
rect 74718 49280 74724 49292
rect 37240 49252 74724 49280
rect 37240 49240 37246 49252
rect 74718 49240 74724 49252
rect 74776 49240 74782 49292
rect 79962 49240 79968 49292
rect 80020 49280 80026 49292
rect 111242 49280 111248 49292
rect 80020 49252 111248 49280
rect 80020 49240 80026 49252
rect 111242 49240 111248 49252
rect 111300 49240 111306 49292
rect 128998 49240 129004 49292
rect 129056 49280 129062 49292
rect 151906 49280 151912 49292
rect 129056 49252 151912 49280
rect 129056 49240 129062 49252
rect 151906 49240 151912 49252
rect 151964 49240 151970 49292
rect 4798 49172 4804 49224
rect 4856 49212 4862 49224
rect 43254 49212 43260 49224
rect 4856 49184 43260 49212
rect 4856 49172 4862 49184
rect 43254 49172 43260 49184
rect 43312 49172 43318 49224
rect 48222 49172 48228 49224
rect 48280 49212 48286 49224
rect 83826 49212 83832 49224
rect 48280 49184 83832 49212
rect 48280 49172 48286 49184
rect 83826 49172 83832 49184
rect 83884 49172 83890 49224
rect 86770 49172 86776 49224
rect 86828 49212 86834 49224
rect 117406 49212 117412 49224
rect 86828 49184 117412 49212
rect 86828 49172 86834 49184
rect 117406 49172 117412 49184
rect 117464 49172 117470 49224
rect 131022 49172 131028 49224
rect 131080 49212 131086 49224
rect 154942 49212 154948 49224
rect 131080 49184 154948 49212
rect 131080 49172 131086 49184
rect 154942 49172 154948 49184
rect 155000 49172 155006 49224
rect 17862 49104 17868 49156
rect 17920 49144 17926 49156
rect 57422 49144 57428 49156
rect 17920 49116 57428 49144
rect 17920 49104 17926 49116
rect 57422 49104 57428 49116
rect 57480 49104 57486 49156
rect 62022 49104 62028 49156
rect 62080 49144 62086 49156
rect 96062 49144 96068 49156
rect 62080 49116 96068 49144
rect 62080 49104 62086 49116
rect 96062 49104 96068 49116
rect 96120 49104 96126 49156
rect 97902 49104 97908 49156
rect 97960 49144 97966 49156
rect 126514 49144 126520 49156
rect 97960 49116 126520 49144
rect 97960 49104 97966 49116
rect 126514 49104 126520 49116
rect 126572 49104 126578 49156
rect 129642 49104 129648 49156
rect 129700 49144 129706 49156
rect 153930 49144 153936 49156
rect 129700 49116 153936 49144
rect 129700 49104 129706 49116
rect 153930 49104 153936 49116
rect 153988 49104 153994 49156
rect 8202 49036 8208 49088
rect 8260 49076 8266 49088
rect 49326 49076 49332 49088
rect 8260 49048 49332 49076
rect 8260 49036 8266 49048
rect 49326 49036 49332 49048
rect 49384 49036 49390 49088
rect 59262 49036 59268 49088
rect 59320 49076 59326 49088
rect 93026 49076 93032 49088
rect 59320 49048 93032 49076
rect 59320 49036 59326 49048
rect 93026 49036 93032 49048
rect 93084 49036 93090 49088
rect 104802 49036 104808 49088
rect 104860 49076 104866 49088
rect 132586 49076 132592 49088
rect 104860 49048 132592 49076
rect 104860 49036 104866 49048
rect 132586 49036 132592 49048
rect 132644 49036 132650 49088
rect 133782 49036 133788 49088
rect 133840 49076 133846 49088
rect 156966 49076 156972 49088
rect 133840 49048 156972 49076
rect 133840 49036 133846 49048
rect 156966 49036 156972 49048
rect 157024 49036 157030 49088
rect 3970 48968 3976 49020
rect 4028 49008 4034 49020
rect 45278 49008 45284 49020
rect 4028 48980 45284 49008
rect 4028 48968 4034 48980
rect 45278 48968 45284 48980
rect 45336 48968 45342 49020
rect 55122 48968 55128 49020
rect 55180 49008 55186 49020
rect 89898 49008 89904 49020
rect 55180 48980 89904 49008
rect 55180 48968 55186 48980
rect 89898 48968 89904 48980
rect 89956 48968 89962 49020
rect 91002 48968 91008 49020
rect 91060 49008 91066 49020
rect 120442 49008 120448 49020
rect 91060 48980 120448 49008
rect 91060 48968 91066 48980
rect 120442 48968 120448 48980
rect 120500 48968 120506 49020
rect 126882 48968 126888 49020
rect 126940 49008 126946 49020
rect 150894 49008 150900 49020
rect 126940 48980 150900 49008
rect 126940 48968 126946 48980
rect 150894 48968 150900 48980
rect 150952 48968 150958 49020
rect 555418 46860 555424 46912
rect 555476 46900 555482 46912
rect 580166 46900 580172 46912
rect 555476 46872 580172 46900
rect 555476 46860 555482 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 293954 46112 293960 46164
rect 294012 46152 294018 46164
rect 294782 46152 294788 46164
rect 294012 46124 294788 46152
rect 294012 46112 294018 46124
rect 294782 46112 294788 46124
rect 294840 46112 294846 46164
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 18598 45540 18604 45552
rect 3476 45512 18604 45540
rect 3476 45500 3482 45512
rect 18598 45500 18604 45512
rect 18656 45500 18662 45552
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 35158 33096 35164 33108
rect 3568 33068 35164 33096
rect 3568 33056 3574 33068
rect 35158 33056 35164 33068
rect 35216 33056 35222 33108
rect 574738 33056 574744 33108
rect 574796 33096 574802 33108
rect 580166 33096 580172 33108
rect 574796 33068 580172 33096
rect 574796 33056 574802 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 108942 22720 108948 22772
rect 109000 22760 109006 22772
rect 134518 22760 134524 22772
rect 109000 22732 134524 22760
rect 109000 22720 109006 22732
rect 134518 22720 134524 22732
rect 134576 22720 134582 22772
rect 30282 21360 30288 21412
rect 30340 21400 30346 21412
rect 67726 21400 67732 21412
rect 30340 21372 67732 21400
rect 30340 21360 30346 21372
rect 67726 21360 67732 21372
rect 67784 21360 67790 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 29638 20652 29644 20664
rect 3476 20624 29644 20652
rect 3476 20612 3482 20624
rect 29638 20612 29644 20624
rect 29696 20612 29702 20664
rect 566458 20612 566464 20664
rect 566516 20652 566522 20664
rect 579982 20652 579988 20664
rect 566516 20624 579988 20652
rect 566516 20612 566522 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 151078 10276 151084 10328
rect 151136 10316 151142 10328
rect 158806 10316 158812 10328
rect 151136 10288 158812 10316
rect 151136 10276 151142 10288
rect 158806 10276 158812 10288
rect 158864 10276 158870 10328
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 21358 6848 21364 6860
rect 3476 6820 21364 6848
rect 3476 6808 3482 6820
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 551278 6808 551284 6860
rect 551336 6848 551342 6860
rect 580166 6848 580172 6860
rect 551336 6820 580172 6848
rect 551336 6808 551342 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 21818 6128 21824 6180
rect 21876 6168 21882 6180
rect 60734 6168 60740 6180
rect 21876 6140 60740 6168
rect 21876 6128 21882 6140
rect 60734 6128 60740 6140
rect 60792 6128 60798 6180
rect 520918 6128 520924 6180
rect 520976 6168 520982 6180
rect 551462 6168 551468 6180
rect 520976 6140 551468 6168
rect 520976 6128 520982 6140
rect 551462 6128 551468 6140
rect 551520 6128 551526 6180
rect 556798 5516 556804 5568
rect 556856 5556 556862 5568
rect 558546 5556 558552 5568
rect 556856 5528 558552 5556
rect 556856 5516 556862 5528
rect 558546 5516 558552 5528
rect 558604 5516 558610 5568
rect 560938 5516 560944 5568
rect 560996 5556 561002 5568
rect 562042 5556 562048 5568
rect 560996 5528 562048 5556
rect 560996 5516 561002 5528
rect 562042 5516 562048 5528
rect 562100 5516 562106 5568
rect 504358 5380 504364 5432
rect 504416 5420 504422 5432
rect 526622 5420 526628 5432
rect 504416 5392 526628 5420
rect 504416 5380 504422 5392
rect 526622 5380 526628 5392
rect 526680 5380 526686 5432
rect 500218 5312 500224 5364
rect 500276 5352 500282 5364
rect 523034 5352 523040 5364
rect 500276 5324 523040 5352
rect 500276 5312 500282 5324
rect 523034 5312 523040 5324
rect 523092 5312 523098 5364
rect 482278 5244 482284 5296
rect 482336 5284 482342 5296
rect 505370 5284 505376 5296
rect 482336 5256 505376 5284
rect 482336 5244 482342 5256
rect 505370 5244 505376 5256
rect 505428 5244 505434 5296
rect 461578 5176 461584 5228
rect 461636 5216 461642 5228
rect 484026 5216 484032 5228
rect 461636 5188 484032 5216
rect 461636 5176 461642 5188
rect 484026 5176 484032 5188
rect 484084 5176 484090 5228
rect 487062 5176 487068 5228
rect 487120 5216 487126 5228
rect 515950 5216 515956 5228
rect 487120 5188 515956 5216
rect 487120 5176 487126 5188
rect 515950 5176 515956 5188
rect 516008 5176 516014 5228
rect 446398 5108 446404 5160
rect 446456 5148 446462 5160
rect 462774 5148 462780 5160
rect 446456 5120 462780 5148
rect 446456 5108 446462 5120
rect 462774 5108 462780 5120
rect 462832 5108 462838 5160
rect 480070 5108 480076 5160
rect 480128 5148 480134 5160
rect 508866 5148 508872 5160
rect 480128 5120 508872 5148
rect 480128 5108 480134 5120
rect 508866 5108 508872 5120
rect 508924 5108 508930 5160
rect 462222 5040 462228 5092
rect 462280 5080 462286 5092
rect 487614 5080 487620 5092
rect 462280 5052 487620 5080
rect 462280 5040 462286 5052
rect 487614 5040 487620 5052
rect 487672 5040 487678 5092
rect 489822 5040 489828 5092
rect 489880 5080 489886 5092
rect 519446 5080 519452 5092
rect 489880 5052 519452 5080
rect 489880 5040 489886 5052
rect 519446 5040 519452 5052
rect 519504 5040 519510 5092
rect 519538 5040 519544 5092
rect 519596 5080 519602 5092
rect 547874 5080 547880 5092
rect 519596 5052 547880 5080
rect 519596 5040 519602 5052
rect 547874 5040 547880 5052
rect 547932 5040 547938 5092
rect 431862 4972 431868 5024
rect 431920 5012 431926 5024
rect 452102 5012 452108 5024
rect 431920 4984 452108 5012
rect 431920 4972 431926 4984
rect 452102 4972 452108 4984
rect 452160 4972 452166 5024
rect 464890 4972 464896 5024
rect 464948 5012 464954 5024
rect 491018 5012 491024 5024
rect 464948 4984 491024 5012
rect 464948 4972 464954 4984
rect 491018 4972 491024 4984
rect 491076 4972 491082 5024
rect 502242 4972 502248 5024
rect 502300 5012 502306 5024
rect 533706 5012 533712 5024
rect 502300 4984 533712 5012
rect 502300 4972 502306 4984
rect 533706 4972 533712 4984
rect 533764 4972 533770 5024
rect 536098 4972 536104 5024
rect 536156 5012 536162 5024
rect 544378 5012 544384 5024
rect 536156 4984 544384 5012
rect 536156 4972 536162 4984
rect 544378 4972 544384 4984
rect 544436 4972 544442 5024
rect 429102 4904 429108 4956
rect 429160 4944 429166 4956
rect 448606 4944 448612 4956
rect 429160 4916 448612 4944
rect 429160 4904 429166 4916
rect 448606 4904 448612 4916
rect 448664 4904 448670 4956
rect 469030 4904 469036 4956
rect 469088 4944 469094 4956
rect 494698 4944 494704 4956
rect 469088 4916 494704 4944
rect 469088 4904 469094 4916
rect 494698 4904 494704 4916
rect 494756 4904 494762 4956
rect 505002 4904 505008 4956
rect 505060 4944 505066 4956
rect 537202 4944 537208 4956
rect 505060 4916 537208 4944
rect 505060 4904 505066 4916
rect 537202 4904 537208 4916
rect 537260 4904 537266 4956
rect 93946 4836 93952 4888
rect 94004 4876 94010 4888
rect 122834 4876 122840 4888
rect 94004 4848 122840 4876
rect 94004 4836 94010 4848
rect 122834 4836 122840 4848
rect 122892 4836 122898 4888
rect 437290 4836 437296 4888
rect 437348 4876 437354 4888
rect 459186 4876 459192 4888
rect 437348 4848 459192 4876
rect 437348 4836 437354 4848
rect 459186 4836 459192 4848
rect 459244 4836 459250 4888
rect 471790 4836 471796 4888
rect 471848 4876 471854 4888
rect 498194 4876 498200 4888
rect 471848 4848 498200 4876
rect 471848 4836 471854 4848
rect 498194 4836 498200 4848
rect 498252 4836 498258 4888
rect 507762 4836 507768 4888
rect 507820 4876 507826 4888
rect 540790 4876 540796 4888
rect 507820 4848 540796 4876
rect 507820 4836 507826 4848
rect 540790 4836 540796 4848
rect 540848 4836 540854 4888
rect 76190 4768 76196 4820
rect 76248 4808 76254 4820
rect 107654 4808 107660 4820
rect 76248 4780 107660 4808
rect 76248 4768 76254 4780
rect 107654 4768 107660 4780
rect 107712 4768 107718 4820
rect 435358 4768 435364 4820
rect 435416 4808 435422 4820
rect 455690 4808 455696 4820
rect 435416 4780 455696 4808
rect 435416 4768 435422 4780
rect 455690 4768 455696 4780
rect 455748 4768 455754 4820
rect 457438 4768 457444 4820
rect 457496 4808 457502 4820
rect 480530 4808 480536 4820
rect 457496 4780 480536 4808
rect 457496 4768 457502 4780
rect 480530 4768 480536 4780
rect 480588 4768 480594 4820
rect 484210 4768 484216 4820
rect 484268 4808 484274 4820
rect 512454 4808 512460 4820
rect 484268 4780 512460 4808
rect 484268 4768 484274 4780
rect 512454 4768 512460 4780
rect 512512 4768 512518 4820
rect 518710 4768 518716 4820
rect 518768 4808 518774 4820
rect 552658 4808 552664 4820
rect 518768 4780 552664 4808
rect 518768 4768 518774 4780
rect 552658 4768 552664 4780
rect 552716 4768 552722 4820
rect 62114 4632 62120 4684
rect 62172 4672 62178 4684
rect 64874 4672 64880 4684
rect 62172 4644 64880 4672
rect 62172 4632 62178 4644
rect 64874 4632 64880 4644
rect 64932 4632 64938 4684
rect 525058 4632 525064 4684
rect 525116 4672 525122 4684
rect 530118 4672 530124 4684
rect 525116 4644 530124 4672
rect 525116 4632 525122 4644
rect 530118 4632 530124 4644
rect 530176 4632 530182 4684
rect 51074 4496 51080 4548
rect 51132 4536 51138 4548
rect 52454 4536 52460 4548
rect 51132 4508 52460 4536
rect 51132 4496 51138 4508
rect 52454 4496 52460 4508
rect 52512 4496 52518 4548
rect 493318 4428 493324 4480
rect 493376 4468 493382 4480
rect 501782 4468 501788 4480
rect 493376 4440 501788 4468
rect 493376 4428 493382 4440
rect 501782 4428 501788 4440
rect 501840 4428 501846 4480
rect 38378 4088 38384 4140
rect 38436 4128 38442 4140
rect 50338 4128 50344 4140
rect 38436 4100 50344 4128
rect 38436 4088 38442 4100
rect 50338 4088 50344 4100
rect 50396 4088 50402 4140
rect 342162 4088 342168 4140
rect 342220 4128 342226 4140
rect 346946 4128 346952 4140
rect 342220 4100 346952 4128
rect 342220 4088 342226 4100
rect 346946 4088 346952 4100
rect 347004 4088 347010 4140
rect 348970 4088 348976 4140
rect 349028 4128 349034 4140
rect 355226 4128 355232 4140
rect 349028 4100 355232 4128
rect 349028 4088 349034 4100
rect 355226 4088 355232 4100
rect 355284 4088 355290 4140
rect 365622 4088 365628 4140
rect 365680 4128 365686 4140
rect 375282 4128 375288 4140
rect 365680 4100 375288 4128
rect 365680 4088 365686 4100
rect 375282 4088 375288 4100
rect 375340 4088 375346 4140
rect 378042 4088 378048 4140
rect 378100 4128 378106 4140
rect 389450 4128 389456 4140
rect 378100 4100 389456 4128
rect 378100 4088 378106 4100
rect 389450 4088 389456 4100
rect 389508 4088 389514 4140
rect 397362 4088 397368 4140
rect 397420 4128 397426 4140
rect 411898 4128 411904 4140
rect 397420 4100 411904 4128
rect 397420 4088 397426 4100
rect 411898 4088 411904 4100
rect 411956 4088 411962 4140
rect 415302 4088 415308 4140
rect 415360 4128 415366 4140
rect 432046 4128 432052 4140
rect 415360 4100 432052 4128
rect 415360 4088 415366 4100
rect 432046 4088 432052 4100
rect 432104 4088 432110 4140
rect 433242 4088 433248 4140
rect 433300 4128 433306 4140
rect 453298 4128 453304 4140
rect 433300 4100 453304 4128
rect 433300 4088 433306 4100
rect 453298 4088 453304 4100
rect 453356 4088 453362 4140
rect 453853 4131 453911 4137
rect 453853 4097 453865 4131
rect 453899 4128 453911 4131
rect 460382 4128 460388 4140
rect 453899 4100 460388 4128
rect 453899 4097 453911 4100
rect 453853 4091 453911 4097
rect 460382 4088 460388 4100
rect 460440 4088 460446 4140
rect 460750 4088 460756 4140
rect 460808 4128 460814 4140
rect 485222 4128 485228 4140
rect 460808 4100 485228 4128
rect 460808 4088 460814 4100
rect 485222 4088 485228 4100
rect 485280 4088 485286 4140
rect 485682 4088 485688 4140
rect 485740 4128 485746 4140
rect 514754 4128 514760 4140
rect 485740 4100 514760 4128
rect 485740 4088 485746 4100
rect 514754 4088 514760 4100
rect 514812 4088 514818 4140
rect 515398 4088 515404 4140
rect 515456 4128 515462 4140
rect 525426 4128 525432 4140
rect 515456 4100 525432 4128
rect 515456 4088 515462 4100
rect 525426 4088 525432 4100
rect 525484 4088 525490 4140
rect 525702 4088 525708 4140
rect 525760 4128 525766 4140
rect 560846 4128 560852 4140
rect 525760 4100 560852 4128
rect 525760 4088 525766 4100
rect 560846 4088 560852 4100
rect 560904 4088 560910 4140
rect 1670 4020 1676 4072
rect 1728 4060 1734 4072
rect 7558 4060 7564 4072
rect 1728 4032 7564 4060
rect 1728 4020 1734 4032
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 41874 4020 41880 4072
rect 41932 4060 41938 4072
rect 50249 4063 50307 4069
rect 50249 4060 50261 4063
rect 41932 4032 50261 4060
rect 41932 4020 41938 4032
rect 50249 4029 50261 4032
rect 50295 4029 50307 4063
rect 50249 4023 50307 4029
rect 53650 4020 53656 4072
rect 53708 4060 53714 4072
rect 64138 4060 64144 4072
rect 53708 4032 64144 4060
rect 53708 4020 53714 4032
rect 64138 4020 64144 4032
rect 64196 4020 64202 4072
rect 314562 4020 314568 4072
rect 314620 4060 314626 4072
rect 316218 4060 316224 4072
rect 314620 4032 316224 4060
rect 314620 4020 314626 4032
rect 316218 4020 316224 4032
rect 316276 4020 316282 4072
rect 332502 4020 332508 4072
rect 332560 4060 332566 4072
rect 336274 4060 336280 4072
rect 332560 4032 336280 4060
rect 332560 4020 332566 4032
rect 336274 4020 336280 4032
rect 336332 4020 336338 4072
rect 340782 4020 340788 4072
rect 340840 4060 340846 4072
rect 345750 4060 345756 4072
rect 340840 4032 345756 4060
rect 340840 4020 340846 4032
rect 345750 4020 345756 4032
rect 345808 4020 345814 4072
rect 351822 4020 351828 4072
rect 351880 4060 351886 4072
rect 358722 4060 358728 4072
rect 351880 4032 358728 4060
rect 351880 4020 351886 4032
rect 358722 4020 358728 4032
rect 358780 4020 358786 4072
rect 367002 4020 367008 4072
rect 367060 4060 367066 4072
rect 376478 4060 376484 4072
rect 367060 4032 376484 4060
rect 367060 4020 367066 4032
rect 376478 4020 376484 4032
rect 376536 4020 376542 4072
rect 382182 4020 382188 4072
rect 382240 4060 382246 4072
rect 394234 4060 394240 4072
rect 382240 4032 394240 4060
rect 382240 4020 382246 4032
rect 394234 4020 394240 4032
rect 394292 4020 394298 4072
rect 395982 4020 395988 4072
rect 396040 4060 396046 4072
rect 410794 4060 410800 4072
rect 396040 4032 410800 4060
rect 396040 4020 396046 4032
rect 410794 4020 410800 4032
rect 410852 4020 410858 4072
rect 411162 4020 411168 4072
rect 411220 4060 411226 4072
rect 428458 4060 428464 4072
rect 411220 4032 428464 4060
rect 411220 4020 411226 4032
rect 428458 4020 428464 4032
rect 428516 4020 428522 4072
rect 430390 4020 430396 4072
rect 430448 4060 430454 4072
rect 450906 4060 450912 4072
rect 430448 4032 450912 4060
rect 430448 4020 430454 4032
rect 450906 4020 450912 4032
rect 450964 4020 450970 4072
rect 456702 4020 456708 4072
rect 456760 4060 456766 4072
rect 481726 4060 481732 4072
rect 456760 4032 481732 4060
rect 456760 4020 456766 4032
rect 481726 4020 481732 4032
rect 481784 4020 481790 4072
rect 484302 4020 484308 4072
rect 484360 4060 484366 4072
rect 513558 4060 513564 4072
rect 484360 4032 513564 4060
rect 484360 4020 484366 4032
rect 513558 4020 513564 4032
rect 513616 4020 513622 4072
rect 518802 4020 518808 4072
rect 518860 4060 518866 4072
rect 548521 4063 548579 4069
rect 548521 4060 548533 4063
rect 518860 4032 548533 4060
rect 518860 4020 518866 4032
rect 548521 4029 548533 4032
rect 548567 4029 548579 4063
rect 548521 4023 548579 4029
rect 548610 4020 548616 4072
rect 548668 4060 548674 4072
rect 549162 4060 549168 4072
rect 548668 4032 549168 4060
rect 548668 4020 548674 4032
rect 549162 4020 549168 4032
rect 549220 4020 549226 4072
rect 31294 3952 31300 4004
rect 31352 3992 31358 4004
rect 43438 3992 43444 4004
rect 31352 3964 43444 3992
rect 31352 3952 31358 3964
rect 43438 3952 43444 3964
rect 43496 3952 43502 4004
rect 45370 3952 45376 4004
rect 45428 3992 45434 4004
rect 71038 3992 71044 4004
rect 45428 3964 71044 3992
rect 45428 3952 45434 3964
rect 71038 3952 71044 3964
rect 71096 3952 71102 4004
rect 92750 3952 92756 4004
rect 92808 3992 92814 4004
rect 95878 3992 95884 4004
rect 92808 3964 95884 3992
rect 92808 3952 92814 3964
rect 95878 3952 95884 3964
rect 95936 3952 95942 4004
rect 357342 3952 357348 4004
rect 357400 3992 357406 4004
rect 364610 3992 364616 4004
rect 357400 3964 364616 3992
rect 357400 3952 357406 3964
rect 364610 3952 364616 3964
rect 364668 3952 364674 4004
rect 372522 3952 372528 4004
rect 372580 3992 372586 4004
rect 382366 3992 382372 4004
rect 372580 3964 382372 3992
rect 372580 3952 372586 3964
rect 382366 3952 382372 3964
rect 382424 3952 382430 4004
rect 383470 3952 383476 4004
rect 383528 3992 383534 4004
rect 395338 3992 395344 4004
rect 383528 3964 395344 3992
rect 383528 3952 383534 3964
rect 395338 3952 395344 3964
rect 395396 3952 395402 4004
rect 398650 3952 398656 4004
rect 398708 3992 398714 4004
rect 413094 3992 413100 4004
rect 398708 3964 413100 3992
rect 398708 3952 398714 3964
rect 413094 3952 413100 3964
rect 413152 3952 413158 4004
rect 415210 3952 415216 4004
rect 415268 3992 415274 4004
rect 433242 3992 433248 4004
rect 415268 3964 433248 3992
rect 415268 3952 415274 3964
rect 433242 3952 433248 3964
rect 433300 3952 433306 4004
rect 436002 3952 436008 4004
rect 436060 3992 436066 4004
rect 456886 3992 456892 4004
rect 436060 3964 456892 3992
rect 436060 3952 436066 3964
rect 456886 3952 456892 3964
rect 456944 3952 456950 4004
rect 463602 3952 463608 4004
rect 463660 3992 463666 4004
rect 488810 3992 488816 4004
rect 463660 3964 488816 3992
rect 463660 3952 463666 3964
rect 488810 3952 488816 3964
rect 488868 3952 488874 4004
rect 493962 3952 493968 4004
rect 494020 3992 494026 4004
rect 524230 3992 524236 4004
rect 494020 3964 524236 3992
rect 494020 3952 494026 3964
rect 524230 3952 524236 3964
rect 524288 3952 524294 4004
rect 524322 3952 524328 4004
rect 524380 3992 524386 4004
rect 559742 3992 559748 4004
rect 524380 3964 559748 3992
rect 524380 3952 524386 3964
rect 559742 3952 559748 3964
rect 559800 3952 559806 4004
rect 28810 3884 28816 3936
rect 28868 3924 28874 3936
rect 55858 3924 55864 3936
rect 28868 3896 55864 3924
rect 28868 3884 28874 3896
rect 55858 3884 55864 3896
rect 55916 3884 55922 3936
rect 71498 3884 71504 3936
rect 71556 3924 71562 3936
rect 75178 3924 75184 3936
rect 71556 3896 75184 3924
rect 71556 3884 71562 3896
rect 75178 3884 75184 3896
rect 75236 3884 75242 3936
rect 353202 3884 353208 3936
rect 353260 3924 353266 3936
rect 361114 3924 361120 3936
rect 353260 3896 361120 3924
rect 353260 3884 353266 3896
rect 361114 3884 361120 3896
rect 361172 3884 361178 3936
rect 362862 3884 362868 3936
rect 362920 3924 362926 3936
rect 371694 3924 371700 3936
rect 362920 3896 371700 3924
rect 362920 3884 362926 3896
rect 371694 3884 371700 3896
rect 371752 3884 371758 3936
rect 373902 3884 373908 3936
rect 373960 3924 373966 3936
rect 384758 3924 384764 3936
rect 373960 3896 384764 3924
rect 373960 3884 373966 3896
rect 384758 3884 384764 3896
rect 384816 3884 384822 3936
rect 384942 3884 384948 3936
rect 385000 3924 385006 3936
rect 397730 3924 397736 3936
rect 385000 3896 397736 3924
rect 385000 3884 385006 3896
rect 397730 3884 397736 3896
rect 397788 3884 397794 3936
rect 400122 3884 400128 3936
rect 400180 3924 400186 3936
rect 415486 3924 415492 3936
rect 400180 3896 415492 3924
rect 400180 3884 400186 3896
rect 415486 3884 415492 3896
rect 415544 3884 415550 3936
rect 419442 3884 419448 3936
rect 419500 3924 419506 3936
rect 437934 3924 437940 3936
rect 419500 3896 437940 3924
rect 419500 3884 419506 3896
rect 437934 3884 437940 3896
rect 437992 3884 437998 3936
rect 438762 3884 438768 3936
rect 438820 3924 438826 3936
rect 453853 3927 453911 3933
rect 453853 3924 453865 3927
rect 438820 3896 453865 3924
rect 438820 3884 438826 3896
rect 453853 3893 453865 3896
rect 453899 3893 453911 3927
rect 453853 3887 453911 3893
rect 453942 3884 453948 3936
rect 454000 3924 454006 3936
rect 458361 3927 458419 3933
rect 458361 3924 458373 3927
rect 454000 3896 458373 3924
rect 454000 3884 454006 3896
rect 458361 3893 458373 3896
rect 458407 3893 458419 3927
rect 458361 3887 458419 3893
rect 460842 3884 460848 3936
rect 460900 3924 460906 3936
rect 486418 3924 486424 3936
rect 460900 3896 486424 3924
rect 460900 3884 460906 3896
rect 486418 3884 486424 3896
rect 486476 3884 486482 3936
rect 491110 3884 491116 3936
rect 491168 3924 491174 3936
rect 520734 3924 520740 3936
rect 491168 3896 520740 3924
rect 491168 3884 491174 3896
rect 520734 3884 520740 3896
rect 520792 3884 520798 3936
rect 521562 3884 521568 3936
rect 521620 3924 521626 3936
rect 548429 3927 548487 3933
rect 548429 3924 548441 3927
rect 521620 3896 548441 3924
rect 521620 3884 521626 3896
rect 548429 3893 548441 3896
rect 548475 3893 548487 3927
rect 548429 3887 548487 3893
rect 548521 3927 548579 3933
rect 548521 3893 548533 3927
rect 548567 3924 548579 3927
rect 553762 3924 553768 3936
rect 548567 3896 553768 3924
rect 548567 3893 548579 3896
rect 548521 3887 548579 3893
rect 553762 3884 553768 3896
rect 553820 3884 553826 3936
rect 24210 3816 24216 3868
rect 24268 3856 24274 3868
rect 54478 3856 54484 3868
rect 24268 3828 54484 3856
rect 24268 3816 24274 3828
rect 54478 3816 54484 3828
rect 54536 3816 54542 3868
rect 353110 3816 353116 3868
rect 353168 3856 353174 3868
rect 359918 3856 359924 3868
rect 353168 3828 359924 3856
rect 353168 3816 353174 3828
rect 359918 3816 359924 3828
rect 359976 3816 359982 3868
rect 360102 3816 360108 3868
rect 360160 3856 360166 3868
rect 368198 3856 368204 3868
rect 360160 3828 368204 3856
rect 360160 3816 360166 3828
rect 368198 3816 368204 3828
rect 368256 3816 368262 3868
rect 371142 3816 371148 3868
rect 371200 3856 371206 3868
rect 381170 3856 381176 3868
rect 371200 3828 381176 3856
rect 371200 3816 371206 3828
rect 381170 3816 381176 3828
rect 381228 3816 381234 3868
rect 386322 3816 386328 3868
rect 386380 3856 386386 3868
rect 398926 3856 398932 3868
rect 386380 3828 398932 3856
rect 386380 3816 386386 3828
rect 398926 3816 398932 3828
rect 398984 3816 398990 3868
rect 405642 3816 405648 3868
rect 405700 3856 405706 3868
rect 421374 3856 421380 3868
rect 405700 3828 421380 3856
rect 405700 3816 405706 3828
rect 421374 3816 421380 3828
rect 421432 3816 421438 3868
rect 424962 3816 424968 3868
rect 425020 3856 425026 3868
rect 443822 3856 443828 3868
rect 425020 3828 443828 3856
rect 425020 3816 425026 3828
rect 443822 3816 443828 3828
rect 443880 3816 443886 3868
rect 448422 3816 448428 3868
rect 448480 3856 448486 3868
rect 471054 3856 471060 3868
rect 448480 3828 471060 3856
rect 448480 3816 448486 3828
rect 471054 3816 471060 3828
rect 471112 3816 471118 3868
rect 471882 3816 471888 3868
rect 471940 3856 471946 3868
rect 499390 3856 499396 3868
rect 471940 3828 499396 3856
rect 471940 3816 471946 3828
rect 499390 3816 499396 3828
rect 499448 3816 499454 3868
rect 500862 3816 500868 3868
rect 500920 3856 500926 3868
rect 532510 3856 532516 3868
rect 500920 3828 532516 3856
rect 500920 3816 500926 3828
rect 532510 3816 532516 3828
rect 532568 3816 532574 3868
rect 538122 3816 538128 3868
rect 538180 3856 538186 3868
rect 575106 3856 575112 3868
rect 538180 3828 575112 3856
rect 538180 3816 538186 3828
rect 575106 3816 575112 3828
rect 575164 3816 575170 3868
rect 20530 3748 20536 3800
rect 20588 3788 20594 3800
rect 44818 3788 44824 3800
rect 20588 3760 44824 3788
rect 20588 3748 20594 3760
rect 44818 3748 44824 3760
rect 44876 3748 44882 3800
rect 46658 3748 46664 3800
rect 46716 3788 46722 3800
rect 76558 3788 76564 3800
rect 46716 3760 76564 3788
rect 46716 3748 46722 3760
rect 76558 3748 76564 3760
rect 76616 3748 76622 3800
rect 344922 3748 344928 3800
rect 344980 3788 344986 3800
rect 351638 3788 351644 3800
rect 344980 3760 351644 3788
rect 344980 3748 344986 3760
rect 351638 3748 351644 3760
rect 351696 3748 351702 3800
rect 358630 3748 358636 3800
rect 358688 3788 358694 3800
rect 367002 3788 367008 3800
rect 358688 3760 367008 3788
rect 358688 3748 358694 3760
rect 367002 3748 367008 3760
rect 367060 3748 367066 3800
rect 368290 3748 368296 3800
rect 368348 3788 368354 3800
rect 377674 3788 377680 3800
rect 368348 3760 377680 3788
rect 368348 3748 368354 3760
rect 377674 3748 377680 3760
rect 377732 3748 377738 3800
rect 380802 3748 380808 3800
rect 380860 3788 380866 3800
rect 393038 3788 393044 3800
rect 380860 3760 393044 3788
rect 380860 3748 380866 3760
rect 393038 3748 393044 3760
rect 393096 3748 393102 3800
rect 393222 3748 393228 3800
rect 393280 3788 393286 3800
rect 407206 3788 407212 3800
rect 393280 3760 407212 3788
rect 393280 3748 393286 3760
rect 407206 3748 407212 3760
rect 407264 3748 407270 3800
rect 411070 3748 411076 3800
rect 411128 3788 411134 3800
rect 427262 3788 427268 3800
rect 411128 3760 427268 3788
rect 411128 3748 411134 3760
rect 427262 3748 427268 3760
rect 427320 3748 427326 3800
rect 427722 3748 427728 3800
rect 427780 3788 427786 3800
rect 447410 3788 447416 3800
rect 427780 3760 447416 3788
rect 427780 3748 427786 3760
rect 447410 3748 447416 3760
rect 447468 3748 447474 3800
rect 449802 3748 449808 3800
rect 449860 3788 449866 3800
rect 472250 3788 472256 3800
rect 449860 3760 472256 3788
rect 449860 3748 449866 3760
rect 472250 3748 472256 3760
rect 472308 3748 472314 3800
rect 475930 3748 475936 3800
rect 475988 3788 475994 3800
rect 502978 3788 502984 3800
rect 475988 3760 502984 3788
rect 475988 3748 475994 3760
rect 502978 3748 502984 3760
rect 503036 3748 503042 3800
rect 503622 3748 503628 3800
rect 503680 3788 503686 3800
rect 534902 3788 534908 3800
rect 503680 3760 534908 3788
rect 503680 3748 503686 3760
rect 534902 3748 534908 3760
rect 534960 3748 534966 3800
rect 536742 3748 536748 3800
rect 536800 3788 536806 3800
rect 573910 3788 573916 3800
rect 536800 3760 573916 3788
rect 536800 3748 536806 3760
rect 573910 3748 573916 3760
rect 573968 3748 573974 3800
rect 35986 3680 35992 3732
rect 36044 3720 36050 3732
rect 71130 3720 71136 3732
rect 36044 3692 71136 3720
rect 36044 3680 36050 3692
rect 71130 3680 71136 3692
rect 71188 3680 71194 3732
rect 350442 3680 350448 3732
rect 350500 3720 350506 3732
rect 357526 3720 357532 3732
rect 350500 3692 357532 3720
rect 350500 3680 350506 3692
rect 357526 3680 357532 3692
rect 357584 3680 357590 3732
rect 361482 3680 361488 3732
rect 361540 3720 361546 3732
rect 369394 3720 369400 3732
rect 361540 3692 369400 3720
rect 361540 3680 361546 3692
rect 369394 3680 369400 3692
rect 369452 3680 369458 3732
rect 369762 3680 369768 3732
rect 369820 3720 369826 3732
rect 379974 3720 379980 3732
rect 369820 3692 379980 3720
rect 369820 3680 369826 3692
rect 379974 3680 379980 3692
rect 380032 3680 380038 3732
rect 389082 3680 389088 3732
rect 389140 3720 389146 3732
rect 402514 3720 402520 3732
rect 389140 3692 402520 3720
rect 389140 3680 389146 3692
rect 402514 3680 402520 3692
rect 402572 3680 402578 3732
rect 404262 3680 404268 3732
rect 404320 3720 404326 3732
rect 420178 3720 420184 3732
rect 404320 3692 420184 3720
rect 404320 3680 404326 3692
rect 420178 3680 420184 3692
rect 420236 3680 420242 3732
rect 422202 3680 422208 3732
rect 422260 3720 422266 3732
rect 440326 3720 440332 3732
rect 422260 3692 440332 3720
rect 422260 3680 422266 3692
rect 440326 3680 440332 3692
rect 440384 3680 440390 3732
rect 442902 3680 442908 3732
rect 442960 3720 442966 3732
rect 465166 3720 465172 3732
rect 442960 3692 465172 3720
rect 442960 3680 442966 3692
rect 465166 3680 465172 3692
rect 465224 3680 465230 3732
rect 467742 3680 467748 3732
rect 467800 3720 467806 3732
rect 493502 3720 493508 3732
rect 467800 3692 493508 3720
rect 467800 3680 467806 3692
rect 493502 3680 493508 3692
rect 493560 3680 493566 3732
rect 496722 3680 496728 3732
rect 496780 3720 496786 3732
rect 527818 3720 527824 3732
rect 496780 3692 527824 3720
rect 496780 3680 496786 3692
rect 527818 3680 527824 3692
rect 527876 3680 527882 3732
rect 533982 3680 533988 3732
rect 534040 3720 534046 3732
rect 570322 3720 570328 3732
rect 534040 3692 570328 3720
rect 534040 3680 534046 3692
rect 570322 3680 570328 3692
rect 570380 3680 570386 3732
rect 26510 3612 26516 3664
rect 26568 3652 26574 3664
rect 26568 3624 35894 3652
rect 26568 3612 26574 3624
rect 566 3544 572 3596
rect 624 3584 630 3596
rect 4798 3584 4804 3596
rect 624 3556 4804 3584
rect 624 3544 630 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12308 3556 12572 3584
rect 12308 3544 12314 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3878 3516 3884 3528
rect 2924 3488 3884 3516
rect 2924 3476 2930 3488
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12342 3516 12348 3528
rect 11204 3488 12348 3516
rect 11204 3476 11210 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 12544 3516 12572 3556
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 16482 3584 16488 3596
rect 15988 3556 16488 3584
rect 15988 3544 15994 3556
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17862 3584 17868 3596
rect 17092 3556 17868 3584
rect 17092 3544 17098 3556
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 19242 3584 19248 3596
rect 18288 3556 19248 3584
rect 18288 3544 18294 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 20622 3584 20628 3596
rect 19484 3556 20628 3584
rect 19484 3544 19490 3556
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 26142 3584 26148 3596
rect 25372 3556 26148 3584
rect 25372 3544 25378 3556
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28902 3584 28908 3596
rect 27764 3556 28908 3584
rect 27764 3544 27770 3556
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 33042 3584 33048 3596
rect 32456 3556 33048 3584
rect 32456 3544 32462 3556
rect 33042 3544 33048 3556
rect 33100 3544 33106 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 34422 3584 34428 3596
rect 33652 3556 34428 3584
rect 33652 3544 33658 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 35866 3584 35894 3624
rect 43070 3612 43076 3664
rect 43128 3652 43134 3664
rect 78858 3652 78864 3664
rect 43128 3624 78864 3652
rect 43128 3612 43134 3624
rect 78858 3612 78864 3624
rect 78916 3612 78922 3664
rect 96246 3612 96252 3664
rect 96304 3652 96310 3664
rect 98638 3652 98644 3664
rect 96304 3624 98644 3652
rect 96304 3612 96310 3624
rect 98638 3612 98644 3624
rect 98696 3612 98702 3664
rect 151078 3652 151084 3664
rect 142126 3624 151084 3652
rect 62114 3584 62120 3596
rect 35866 3556 62120 3584
rect 62114 3544 62120 3556
rect 62172 3544 62178 3596
rect 66714 3544 66720 3596
rect 66772 3584 66778 3596
rect 67542 3584 67548 3596
rect 66772 3556 67548 3584
rect 66772 3544 66778 3556
rect 67542 3544 67548 3556
rect 67600 3544 67606 3596
rect 67910 3544 67916 3596
rect 67968 3584 67974 3596
rect 68922 3584 68928 3596
rect 67968 3556 68928 3584
rect 67968 3544 67974 3556
rect 68922 3544 68928 3556
rect 68980 3544 68986 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 70210 3584 70216 3596
rect 69164 3556 70216 3584
rect 69164 3544 69170 3556
rect 70210 3544 70216 3556
rect 70268 3544 70274 3596
rect 72602 3544 72608 3596
rect 72660 3584 72666 3596
rect 73062 3584 73068 3596
rect 72660 3556 73068 3584
rect 72660 3544 72666 3556
rect 73062 3544 73068 3556
rect 73120 3544 73126 3596
rect 73798 3544 73804 3596
rect 73856 3584 73862 3596
rect 74442 3584 74448 3596
rect 73856 3556 74448 3584
rect 73856 3544 73862 3556
rect 74442 3544 74448 3556
rect 74500 3544 74506 3596
rect 74994 3544 75000 3596
rect 75052 3584 75058 3596
rect 75822 3584 75828 3596
rect 75052 3556 75828 3584
rect 75052 3544 75058 3556
rect 75822 3544 75828 3556
rect 75880 3544 75886 3596
rect 77386 3544 77392 3596
rect 77444 3584 77450 3596
rect 78582 3584 78588 3596
rect 77444 3556 78588 3584
rect 77444 3544 77450 3556
rect 78582 3544 78588 3556
rect 78640 3544 78646 3596
rect 80882 3544 80888 3596
rect 80940 3584 80946 3596
rect 81342 3584 81348 3596
rect 80940 3556 81348 3584
rect 80940 3544 80946 3556
rect 81342 3544 81348 3556
rect 81400 3544 81406 3596
rect 83274 3544 83280 3596
rect 83332 3584 83338 3596
rect 84102 3584 84108 3596
rect 83332 3556 84108 3584
rect 83332 3544 83338 3556
rect 84102 3544 84108 3556
rect 84160 3544 84166 3596
rect 85666 3544 85672 3596
rect 85724 3584 85730 3596
rect 86770 3584 86776 3596
rect 85724 3556 86776 3584
rect 85724 3544 85730 3556
rect 86770 3544 86776 3556
rect 86828 3544 86834 3596
rect 114002 3544 114008 3596
rect 114060 3584 114066 3596
rect 124858 3584 124864 3596
rect 114060 3556 124864 3584
rect 114060 3544 114066 3556
rect 124858 3544 124864 3556
rect 124916 3544 124922 3596
rect 136450 3544 136456 3596
rect 136508 3584 136514 3596
rect 142126 3584 142154 3624
rect 151078 3612 151084 3624
rect 151136 3612 151142 3664
rect 343542 3612 343548 3664
rect 343600 3652 343606 3664
rect 349246 3652 349252 3664
rect 343600 3624 349252 3652
rect 343600 3612 343606 3624
rect 349246 3612 349252 3624
rect 349304 3612 349310 3664
rect 357250 3612 357256 3664
rect 357308 3652 357314 3664
rect 365806 3652 365812 3664
rect 357308 3624 365812 3652
rect 357308 3612 357314 3624
rect 365806 3612 365812 3624
rect 365864 3612 365870 3664
rect 368382 3612 368388 3664
rect 368440 3652 368446 3664
rect 378870 3652 378876 3664
rect 368440 3624 378876 3652
rect 368440 3612 368446 3624
rect 378870 3612 378876 3624
rect 378928 3612 378934 3664
rect 379422 3612 379428 3664
rect 379480 3652 379486 3664
rect 390646 3652 390652 3664
rect 379480 3624 390652 3652
rect 379480 3612 379486 3624
rect 390646 3612 390652 3624
rect 390704 3612 390710 3664
rect 391750 3612 391756 3664
rect 391808 3652 391814 3664
rect 404814 3652 404820 3664
rect 391808 3624 404820 3652
rect 391808 3612 391814 3624
rect 404814 3612 404820 3624
rect 404872 3612 404878 3664
rect 406930 3612 406936 3664
rect 406988 3652 406994 3664
rect 422570 3652 422576 3664
rect 406988 3624 422576 3652
rect 406988 3612 406994 3624
rect 422570 3612 422576 3624
rect 422628 3612 422634 3664
rect 426250 3612 426256 3664
rect 426308 3652 426314 3664
rect 445018 3652 445024 3664
rect 426308 3624 445024 3652
rect 426308 3612 426314 3624
rect 445018 3612 445024 3624
rect 445076 3612 445082 3664
rect 447042 3612 447048 3664
rect 447100 3652 447106 3664
rect 469858 3652 469864 3664
rect 447100 3624 469864 3652
rect 447100 3612 447106 3624
rect 469858 3612 469864 3624
rect 469916 3612 469922 3664
rect 470502 3612 470508 3664
rect 470560 3652 470566 3664
rect 497090 3652 497096 3664
rect 470560 3624 497096 3652
rect 470560 3612 470566 3624
rect 497090 3612 497096 3624
rect 497148 3612 497154 3664
rect 498102 3612 498108 3664
rect 498160 3652 498166 3664
rect 529014 3652 529020 3664
rect 498160 3624 529020 3652
rect 498160 3612 498166 3624
rect 529014 3612 529020 3624
rect 529072 3612 529078 3664
rect 529842 3612 529848 3664
rect 529900 3652 529906 3664
rect 566826 3652 566832 3664
rect 529900 3624 566832 3652
rect 529900 3612 529906 3624
rect 566826 3612 566832 3624
rect 566884 3612 566890 3664
rect 146938 3584 146944 3596
rect 136508 3556 142154 3584
rect 142356 3556 146944 3584
rect 136508 3544 136514 3556
rect 12544 3488 48912 3516
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 46198 3448 46204 3460
rect 5316 3420 46204 3448
rect 5316 3408 5322 3420
rect 46198 3408 46204 3420
rect 46256 3408 46262 3460
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 44266 3340 44272 3392
rect 44324 3380 44330 3392
rect 45462 3380 45468 3392
rect 44324 3352 45468 3380
rect 44324 3340 44330 3352
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 48884 3380 48912 3488
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 52362 3516 52368 3528
rect 51408 3488 52368 3516
rect 51408 3476 51414 3488
rect 52362 3476 52368 3488
rect 52420 3476 52426 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 53742 3516 53748 3528
rect 52604 3488 53748 3516
rect 52604 3476 52610 3488
rect 53742 3476 53748 3488
rect 53800 3476 53806 3528
rect 57146 3516 57152 3528
rect 55186 3488 57152 3516
rect 50249 3451 50307 3457
rect 50249 3417 50261 3451
rect 50295 3448 50307 3451
rect 55186 3448 55214 3488
rect 57146 3476 57152 3488
rect 57204 3476 57210 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 60826 3476 60832 3528
rect 60884 3516 60890 3528
rect 60884 3488 84424 3516
rect 60884 3476 60890 3488
rect 50295 3420 55214 3448
rect 50295 3417 50307 3420
rect 50249 3411 50307 3417
rect 56042 3408 56048 3460
rect 56100 3448 56106 3460
rect 56502 3448 56508 3460
rect 56100 3420 56508 3448
rect 56100 3408 56106 3420
rect 56502 3408 56508 3420
rect 56560 3408 56566 3460
rect 64322 3408 64328 3460
rect 64380 3448 64386 3460
rect 84396 3448 84424 3488
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 85482 3516 85488 3528
rect 84528 3488 85488 3516
rect 84528 3476 84534 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 90266 3516 90272 3528
rect 89220 3488 90272 3516
rect 89220 3476 89226 3488
rect 90266 3476 90272 3488
rect 90324 3476 90330 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 92382 3516 92388 3528
rect 91612 3488 92388 3516
rect 91612 3476 91618 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 102042 3516 102048 3528
rect 101088 3488 102048 3516
rect 101088 3476 101094 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 102226 3476 102232 3528
rect 102284 3516 102290 3528
rect 103422 3516 103428 3528
rect 102284 3488 103428 3516
rect 102284 3476 102290 3488
rect 103422 3476 103428 3488
rect 103480 3476 103486 3528
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 106182 3516 106188 3528
rect 105780 3488 106188 3516
rect 105780 3476 105786 3488
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 110322 3516 110328 3528
rect 109368 3488 110328 3516
rect 109368 3476 109374 3488
rect 110322 3476 110328 3488
rect 110380 3476 110386 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111702 3516 111708 3528
rect 110564 3488 111708 3516
rect 110564 3476 110570 3488
rect 111702 3476 111708 3488
rect 111760 3476 111766 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 116394 3476 116400 3528
rect 116452 3516 116458 3528
rect 117222 3516 117228 3528
rect 116452 3488 117228 3516
rect 116452 3476 116458 3488
rect 117222 3476 117228 3488
rect 117280 3476 117286 3528
rect 117590 3476 117596 3528
rect 117648 3516 117654 3528
rect 118602 3516 118608 3528
rect 117648 3488 118608 3516
rect 117648 3476 117654 3488
rect 118602 3476 118608 3488
rect 118660 3476 118666 3528
rect 118786 3476 118792 3528
rect 118844 3516 118850 3528
rect 119798 3516 119804 3528
rect 118844 3488 119804 3516
rect 118844 3476 118850 3488
rect 119798 3476 119804 3488
rect 119856 3476 119862 3528
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126882 3516 126888 3528
rect 125928 3488 126888 3516
rect 125928 3476 125934 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128998 3516 129004 3528
rect 127032 3488 129004 3516
rect 127032 3476 127038 3488
rect 128998 3476 129004 3488
rect 129056 3476 129062 3528
rect 130562 3476 130568 3528
rect 130620 3516 130626 3528
rect 131022 3516 131028 3528
rect 130620 3488 131028 3516
rect 130620 3476 130626 3488
rect 131022 3476 131028 3488
rect 131080 3476 131086 3528
rect 142356 3516 142384 3556
rect 146938 3544 146944 3556
rect 146996 3544 147002 3596
rect 267734 3544 267740 3596
rect 267792 3584 267798 3596
rect 268930 3584 268936 3596
rect 267792 3556 268936 3584
rect 267792 3544 267798 3556
rect 268930 3544 268936 3556
rect 268988 3544 268994 3596
rect 324222 3544 324228 3596
rect 324280 3584 324286 3596
rect 326798 3584 326804 3596
rect 324280 3556 326804 3584
rect 324280 3544 324286 3556
rect 326798 3544 326804 3556
rect 326856 3544 326862 3596
rect 328362 3544 328368 3596
rect 328420 3584 328426 3596
rect 331582 3584 331588 3596
rect 328420 3556 331588 3584
rect 328420 3544 328426 3556
rect 331582 3544 331588 3556
rect 331640 3544 331646 3596
rect 334618 3544 334624 3596
rect 334676 3584 334682 3596
rect 338666 3584 338672 3596
rect 334676 3556 338672 3584
rect 334676 3544 334682 3556
rect 338666 3544 338672 3556
rect 338724 3544 338730 3596
rect 339402 3544 339408 3596
rect 339460 3584 339466 3596
rect 344554 3584 344560 3596
rect 339460 3556 344560 3584
rect 339460 3544 339466 3556
rect 344554 3544 344560 3556
rect 344612 3544 344618 3596
rect 354582 3544 354588 3596
rect 354640 3584 354646 3596
rect 362310 3584 362316 3596
rect 354640 3556 362316 3584
rect 354640 3544 354646 3556
rect 362310 3544 362316 3556
rect 362368 3544 362374 3596
rect 364150 3544 364156 3596
rect 364208 3584 364214 3596
rect 372890 3584 372896 3596
rect 364208 3556 372896 3584
rect 364208 3544 364214 3556
rect 372890 3544 372896 3556
rect 372948 3544 372954 3596
rect 376570 3544 376576 3596
rect 376628 3584 376634 3596
rect 387150 3584 387156 3596
rect 376628 3556 387156 3584
rect 376628 3544 376634 3556
rect 387150 3544 387156 3556
rect 387208 3544 387214 3596
rect 387610 3544 387616 3596
rect 387668 3584 387674 3596
rect 401318 3584 401324 3596
rect 387668 3556 401324 3584
rect 387668 3544 387674 3556
rect 401318 3544 401324 3556
rect 401376 3544 401382 3596
rect 402790 3544 402796 3596
rect 402848 3584 402854 3596
rect 418982 3584 418988 3596
rect 402848 3556 418988 3584
rect 402848 3544 402854 3556
rect 418982 3544 418988 3556
rect 419040 3544 419046 3596
rect 422110 3544 422116 3596
rect 422168 3584 422174 3596
rect 441522 3584 441528 3596
rect 422168 3556 441528 3584
rect 422168 3544 422174 3556
rect 441522 3544 441528 3556
rect 441580 3544 441586 3596
rect 441614 3544 441620 3596
rect 441672 3584 441678 3596
rect 463970 3584 463976 3596
rect 441672 3556 463976 3584
rect 441672 3544 441678 3556
rect 463970 3544 463976 3556
rect 464028 3544 464034 3596
rect 464982 3544 464988 3596
rect 465040 3584 465046 3596
rect 489914 3584 489920 3596
rect 465040 3556 489920 3584
rect 465040 3544 465046 3556
rect 489914 3544 489920 3556
rect 489972 3544 489978 3596
rect 491202 3544 491208 3596
rect 491260 3584 491266 3596
rect 521838 3584 521844 3596
rect 491260 3556 521844 3584
rect 491260 3544 491266 3556
rect 521838 3544 521844 3556
rect 521896 3544 521902 3596
rect 527082 3544 527088 3596
rect 527140 3584 527146 3596
rect 563238 3584 563244 3596
rect 527140 3556 563244 3584
rect 527140 3544 527146 3556
rect 563238 3544 563244 3556
rect 563296 3544 563302 3596
rect 132466 3488 142384 3516
rect 88978 3448 88984 3460
rect 64380 3420 84194 3448
rect 84396 3420 88984 3448
rect 64380 3408 64386 3420
rect 51074 3380 51080 3392
rect 48884 3352 51080 3380
rect 51074 3340 51080 3352
rect 51132 3340 51138 3392
rect 78582 3340 78588 3392
rect 78640 3380 78646 3392
rect 81986 3380 81992 3392
rect 78640 3352 81992 3380
rect 78640 3340 78646 3352
rect 81986 3340 81992 3352
rect 82044 3340 82050 3392
rect 82078 3340 82084 3392
rect 82136 3380 82142 3392
rect 83458 3380 83464 3392
rect 82136 3352 83464 3380
rect 82136 3340 82142 3352
rect 83458 3340 83464 3352
rect 83516 3340 83522 3392
rect 84166 3380 84194 3420
rect 88978 3408 88984 3420
rect 89036 3408 89042 3460
rect 103330 3408 103336 3460
rect 103388 3448 103394 3460
rect 106826 3448 106832 3460
rect 103388 3420 106832 3448
rect 103388 3408 103394 3420
rect 106826 3408 106832 3420
rect 106884 3408 106890 3460
rect 111610 3408 111616 3460
rect 111668 3448 111674 3460
rect 111668 3420 122834 3448
rect 111668 3408 111674 3420
rect 93118 3380 93124 3392
rect 84166 3352 93124 3380
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 122806 3380 122834 3420
rect 128170 3408 128176 3460
rect 128228 3448 128234 3460
rect 132466 3448 132494 3488
rect 142430 3476 142436 3528
rect 142488 3516 142494 3528
rect 143442 3516 143448 3528
rect 142488 3488 143448 3516
rect 142488 3476 142494 3488
rect 143442 3476 143448 3488
rect 143500 3476 143506 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144638 3516 144644 3528
rect 143592 3488 144644 3516
rect 143592 3476 143598 3488
rect 144638 3476 144644 3488
rect 144696 3476 144702 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
rect 150342 3516 150348 3528
rect 149572 3488 150348 3516
rect 149572 3476 149578 3488
rect 150342 3476 150348 3488
rect 150400 3476 150406 3528
rect 150618 3476 150624 3528
rect 150676 3516 150682 3528
rect 151722 3516 151728 3528
rect 150676 3488 151728 3516
rect 150676 3476 150682 3488
rect 151722 3476 151728 3488
rect 151780 3476 151786 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 153102 3516 153108 3528
rect 151872 3488 153108 3516
rect 151872 3476 151878 3488
rect 153102 3476 153108 3488
rect 153160 3476 153166 3528
rect 155402 3476 155408 3528
rect 155460 3516 155466 3528
rect 155862 3516 155868 3528
rect 155460 3488 155868 3516
rect 155460 3476 155466 3488
rect 155862 3476 155868 3488
rect 155920 3476 155926 3528
rect 156598 3476 156604 3528
rect 156656 3516 156662 3528
rect 157242 3516 157248 3528
rect 156656 3488 157248 3516
rect 156656 3476 156662 3488
rect 157242 3476 157248 3488
rect 157300 3476 157306 3528
rect 157794 3476 157800 3528
rect 157852 3516 157858 3528
rect 158622 3516 158628 3528
rect 157852 3488 158628 3516
rect 157852 3476 157858 3488
rect 158622 3476 158628 3488
rect 158680 3476 158686 3528
rect 158898 3476 158904 3528
rect 158956 3516 158962 3528
rect 160002 3516 160008 3528
rect 158956 3488 160008 3516
rect 158956 3476 158962 3488
rect 160002 3476 160008 3488
rect 160060 3476 160066 3528
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161382 3516 161388 3528
rect 160152 3488 161388 3516
rect 160152 3476 160158 3488
rect 161382 3476 161388 3488
rect 161440 3476 161446 3528
rect 163682 3476 163688 3528
rect 163740 3516 163746 3528
rect 164142 3516 164148 3528
rect 163740 3488 164148 3516
rect 163740 3476 163746 3488
rect 164142 3476 164148 3488
rect 164200 3476 164206 3528
rect 166074 3476 166080 3528
rect 166132 3516 166138 3528
rect 166902 3516 166908 3528
rect 166132 3488 166908 3516
rect 166132 3476 166138 3488
rect 166902 3476 166908 3488
rect 166960 3476 166966 3528
rect 167178 3476 167184 3528
rect 167236 3516 167242 3528
rect 168282 3516 168288 3528
rect 167236 3488 168288 3516
rect 167236 3476 167242 3488
rect 168282 3476 168288 3488
rect 168340 3476 168346 3528
rect 168374 3476 168380 3528
rect 168432 3516 168438 3528
rect 169478 3516 169484 3528
rect 168432 3488 169484 3516
rect 168432 3476 168438 3488
rect 169478 3476 169484 3488
rect 169536 3476 169542 3528
rect 171962 3476 171968 3528
rect 172020 3516 172026 3528
rect 172422 3516 172428 3528
rect 172020 3488 172428 3516
rect 172020 3476 172026 3488
rect 172422 3476 172428 3488
rect 172480 3476 172486 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173802 3516 173808 3528
rect 173216 3488 173808 3516
rect 173216 3476 173222 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 174262 3476 174268 3528
rect 174320 3516 174326 3528
rect 175182 3516 175188 3528
rect 174320 3488 175188 3516
rect 174320 3476 174326 3488
rect 175182 3476 175188 3488
rect 175240 3476 175246 3528
rect 175458 3476 175464 3528
rect 175516 3516 175522 3528
rect 176562 3516 176568 3528
rect 175516 3488 176568 3516
rect 175516 3476 175522 3488
rect 176562 3476 176568 3488
rect 176620 3476 176626 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177758 3516 177764 3528
rect 176712 3488 177764 3516
rect 176712 3476 176718 3488
rect 177758 3476 177764 3488
rect 177816 3476 177822 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180702 3516 180708 3528
rect 180300 3488 180708 3516
rect 180300 3476 180306 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 181438 3476 181444 3528
rect 181496 3516 181502 3528
rect 182082 3516 182088 3528
rect 181496 3488 182088 3516
rect 181496 3476 181502 3488
rect 182082 3476 182088 3488
rect 182140 3476 182146 3528
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 184934 3476 184940 3528
rect 184992 3516 184998 3528
rect 186222 3516 186228 3528
rect 184992 3488 186228 3516
rect 184992 3476 184998 3488
rect 186222 3476 186228 3488
rect 186280 3476 186286 3528
rect 188522 3476 188528 3528
rect 188580 3516 188586 3528
rect 188982 3516 188988 3528
rect 188580 3488 188988 3516
rect 188580 3476 188586 3488
rect 188982 3476 188988 3488
rect 189040 3476 189046 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 191742 3516 191748 3528
rect 190880 3488 191748 3516
rect 190880 3476 190886 3488
rect 191742 3476 191748 3488
rect 191800 3476 191806 3528
rect 192018 3476 192024 3528
rect 192076 3516 192082 3528
rect 193122 3516 193128 3528
rect 192076 3488 193128 3516
rect 192076 3476 192082 3488
rect 193122 3476 193128 3488
rect 193180 3476 193186 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194318 3516 194324 3528
rect 193272 3488 194324 3516
rect 193272 3476 193278 3488
rect 194318 3476 194324 3488
rect 194376 3476 194382 3528
rect 197906 3476 197912 3528
rect 197964 3516 197970 3528
rect 198642 3516 198648 3528
rect 197964 3488 198648 3516
rect 197964 3476 197970 3488
rect 198642 3476 198648 3488
rect 198700 3476 198706 3528
rect 199102 3476 199108 3528
rect 199160 3516 199166 3528
rect 200022 3516 200028 3528
rect 199160 3488 200028 3516
rect 199160 3476 199166 3488
rect 200022 3476 200028 3488
rect 200080 3476 200086 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 205542 3516 205548 3528
rect 205140 3488 205548 3516
rect 205140 3476 205146 3488
rect 205542 3476 205548 3488
rect 205600 3476 205606 3528
rect 206186 3476 206192 3528
rect 206244 3516 206250 3528
rect 206922 3516 206928 3528
rect 206244 3488 206928 3516
rect 206244 3476 206250 3488
rect 206922 3476 206928 3488
rect 206980 3476 206986 3528
rect 207382 3476 207388 3528
rect 207440 3516 207446 3528
rect 208302 3516 208308 3528
rect 207440 3488 208308 3516
rect 207440 3476 207446 3488
rect 208302 3476 208308 3488
rect 208360 3476 208366 3528
rect 209774 3476 209780 3528
rect 209832 3516 209838 3528
rect 211062 3516 211068 3528
rect 209832 3488 211068 3516
rect 209832 3476 209838 3488
rect 211062 3476 211068 3488
rect 211120 3476 211126 3528
rect 213362 3476 213368 3528
rect 213420 3516 213426 3528
rect 213822 3516 213828 3528
rect 213420 3488 213828 3516
rect 213420 3476 213426 3488
rect 213822 3476 213828 3488
rect 213880 3476 213886 3528
rect 214466 3476 214472 3528
rect 214524 3516 214530 3528
rect 215202 3516 215208 3528
rect 214524 3488 215208 3516
rect 214524 3476 214530 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 216582 3516 216588 3528
rect 215720 3488 216588 3516
rect 215720 3476 215726 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 216858 3476 216864 3528
rect 216916 3516 216922 3528
rect 217962 3516 217968 3528
rect 216916 3488 217968 3516
rect 216916 3476 216922 3488
rect 217962 3476 217968 3488
rect 218020 3476 218026 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 219158 3516 219164 3528
rect 218112 3488 219164 3516
rect 218112 3476 218118 3488
rect 219158 3476 219164 3488
rect 219216 3476 219222 3528
rect 222746 3476 222752 3528
rect 222804 3516 222810 3528
rect 223482 3516 223488 3528
rect 222804 3488 223488 3516
rect 222804 3476 222810 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 224862 3516 224868 3528
rect 224000 3488 224868 3516
rect 224000 3476 224006 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 227622 3516 227628 3528
rect 226392 3488 227628 3516
rect 226392 3476 226398 3488
rect 227622 3476 227628 3488
rect 227680 3476 227686 3528
rect 229830 3476 229836 3528
rect 229888 3516 229894 3528
rect 230382 3516 230388 3528
rect 229888 3488 230388 3516
rect 229888 3476 229894 3488
rect 230382 3476 230388 3488
rect 230440 3476 230446 3528
rect 231026 3476 231032 3528
rect 231084 3516 231090 3528
rect 231762 3516 231768 3528
rect 231084 3488 231768 3516
rect 231084 3476 231090 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 234614 3476 234620 3528
rect 234672 3516 234678 3528
rect 235902 3516 235908 3528
rect 234672 3488 235908 3516
rect 234672 3476 234678 3488
rect 235902 3476 235908 3488
rect 235960 3476 235966 3528
rect 238110 3476 238116 3528
rect 238168 3516 238174 3528
rect 238662 3516 238668 3528
rect 238168 3488 238668 3516
rect 238168 3476 238174 3488
rect 238662 3476 238668 3488
rect 238720 3476 238726 3528
rect 239306 3476 239312 3528
rect 239364 3516 239370 3528
rect 240042 3516 240048 3528
rect 239364 3488 240048 3516
rect 239364 3476 239370 3488
rect 240042 3476 240048 3488
rect 240100 3476 240106 3528
rect 240502 3476 240508 3528
rect 240560 3516 240566 3528
rect 241422 3516 241428 3528
rect 240560 3488 241428 3516
rect 240560 3476 240566 3488
rect 241422 3476 241428 3488
rect 241480 3476 241486 3528
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 243998 3516 244004 3528
rect 242952 3488 244004 3516
rect 242952 3476 242958 3488
rect 243998 3476 244004 3488
rect 244056 3476 244062 3528
rect 247586 3476 247592 3528
rect 247644 3516 247650 3528
rect 248322 3516 248328 3528
rect 247644 3488 248328 3516
rect 247644 3476 247650 3488
rect 248322 3476 248328 3488
rect 248380 3476 248386 3528
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 251082 3516 251088 3528
rect 250036 3488 251088 3516
rect 250036 3476 250042 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 251174 3476 251180 3528
rect 251232 3516 251238 3528
rect 252462 3516 252468 3528
rect 251232 3488 252468 3516
rect 251232 3476 251238 3488
rect 252462 3476 252468 3488
rect 252520 3476 252526 3528
rect 254670 3476 254676 3528
rect 254728 3516 254734 3528
rect 255222 3516 255228 3528
rect 254728 3488 255228 3516
rect 254728 3476 254734 3488
rect 255222 3476 255228 3488
rect 255280 3476 255286 3528
rect 255866 3476 255872 3528
rect 255924 3516 255930 3528
rect 256602 3516 256608 3528
rect 255924 3488 256608 3516
rect 255924 3476 255930 3488
rect 256602 3476 256608 3488
rect 256660 3476 256666 3528
rect 257062 3476 257068 3528
rect 257120 3516 257126 3528
rect 257982 3516 257988 3528
rect 257120 3488 257988 3516
rect 257120 3476 257126 3488
rect 257982 3476 257988 3488
rect 258040 3476 258046 3528
rect 258258 3476 258264 3528
rect 258316 3516 258322 3528
rect 259362 3516 259368 3528
rect 258316 3488 259368 3516
rect 258316 3476 258322 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 259454 3476 259460 3528
rect 259512 3516 259518 3528
rect 260742 3516 260748 3528
rect 259512 3488 260748 3516
rect 259512 3476 259518 3488
rect 260742 3476 260748 3488
rect 260800 3476 260806 3528
rect 262950 3476 262956 3528
rect 263008 3516 263014 3528
rect 263502 3516 263508 3528
rect 263008 3488 263508 3516
rect 263008 3476 263014 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 264882 3516 264888 3528
rect 264204 3488 264888 3516
rect 264204 3476 264210 3488
rect 264882 3476 264888 3488
rect 264940 3476 264946 3528
rect 266538 3476 266544 3528
rect 266596 3516 266602 3528
rect 267642 3516 267648 3528
rect 266596 3488 267648 3516
rect 266596 3476 266602 3488
rect 267642 3476 267648 3488
rect 267700 3476 267706 3528
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 274542 3516 274548 3528
rect 273680 3488 274548 3516
rect 273680 3476 273686 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 274818 3476 274824 3528
rect 274876 3516 274882 3528
rect 275922 3516 275928 3528
rect 274876 3488 275928 3516
rect 274876 3476 274882 3488
rect 275922 3476 275928 3488
rect 275980 3476 275986 3528
rect 280706 3476 280712 3528
rect 280764 3516 280770 3528
rect 281442 3516 281448 3528
rect 280764 3488 281448 3516
rect 280764 3476 280770 3488
rect 281442 3476 281448 3488
rect 281500 3476 281506 3528
rect 281902 3476 281908 3528
rect 281960 3516 281966 3528
rect 282822 3516 282828 3528
rect 281960 3488 282828 3516
rect 281960 3476 281966 3488
rect 282822 3476 282828 3488
rect 282880 3476 282886 3528
rect 284294 3476 284300 3528
rect 284352 3516 284358 3528
rect 285582 3516 285588 3528
rect 284352 3488 285588 3516
rect 284352 3476 284358 3488
rect 285582 3476 285588 3488
rect 285640 3476 285646 3528
rect 287790 3476 287796 3528
rect 287848 3516 287854 3528
rect 288342 3516 288348 3528
rect 287848 3488 288348 3516
rect 287848 3476 287854 3488
rect 288342 3476 288348 3488
rect 288400 3476 288406 3528
rect 288986 3476 288992 3528
rect 289044 3516 289050 3528
rect 289722 3516 289728 3528
rect 289044 3488 289728 3516
rect 289044 3476 289050 3488
rect 289722 3476 289728 3488
rect 289780 3476 289786 3528
rect 290182 3476 290188 3528
rect 290240 3516 290246 3528
rect 291286 3516 291292 3528
rect 290240 3488 291292 3516
rect 290240 3476 290246 3488
rect 291286 3476 291292 3488
rect 291344 3476 291350 3528
rect 291378 3476 291384 3528
rect 291436 3516 291442 3528
rect 292482 3516 292488 3528
rect 291436 3488 292488 3516
rect 291436 3476 291442 3488
rect 292482 3476 292488 3488
rect 292540 3476 292546 3528
rect 292574 3476 292580 3528
rect 292632 3516 292638 3528
rect 294046 3516 294052 3528
rect 292632 3488 294052 3516
rect 292632 3476 292638 3488
rect 294046 3476 294052 3488
rect 294104 3476 294110 3528
rect 296070 3476 296076 3528
rect 296128 3516 296134 3528
rect 296622 3516 296628 3528
rect 296128 3488 296628 3516
rect 296128 3476 296134 3488
rect 296622 3476 296628 3488
rect 296680 3476 296686 3528
rect 302418 3476 302424 3528
rect 302476 3516 302482 3528
rect 303154 3516 303160 3528
rect 302476 3488 303160 3516
rect 302476 3476 302482 3488
rect 303154 3476 303160 3488
rect 303212 3476 303218 3528
rect 307754 3476 307760 3528
rect 307812 3516 307818 3528
rect 309042 3516 309048 3528
rect 307812 3488 309048 3516
rect 307812 3476 307818 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 310422 3476 310428 3528
rect 310480 3516 310486 3528
rect 311434 3516 311440 3528
rect 310480 3488 311440 3516
rect 310480 3476 310486 3488
rect 311434 3476 311440 3488
rect 311492 3476 311498 3528
rect 311802 3476 311808 3528
rect 311860 3516 311866 3528
rect 312630 3516 312636 3528
rect 311860 3488 312636 3516
rect 311860 3476 311866 3488
rect 312630 3476 312636 3488
rect 312688 3476 312694 3528
rect 314470 3476 314476 3528
rect 314528 3516 314534 3528
rect 315022 3516 315028 3528
rect 314528 3488 315028 3516
rect 314528 3476 314534 3488
rect 315022 3476 315028 3488
rect 315080 3476 315086 3528
rect 318702 3476 318708 3528
rect 318760 3516 318766 3528
rect 319714 3516 319720 3528
rect 318760 3488 319720 3516
rect 318760 3476 318766 3488
rect 319714 3476 319720 3488
rect 319772 3476 319778 3528
rect 322750 3476 322756 3528
rect 322808 3516 322814 3528
rect 324406 3516 324412 3528
rect 322808 3488 324412 3516
rect 322808 3476 322814 3488
rect 324406 3476 324412 3488
rect 324464 3476 324470 3528
rect 329742 3476 329748 3528
rect 329800 3516 329806 3528
rect 332686 3516 332692 3528
rect 329800 3488 332692 3516
rect 329800 3476 329806 3488
rect 332686 3476 332692 3488
rect 332744 3476 332750 3528
rect 335262 3476 335268 3528
rect 335320 3516 335326 3528
rect 335320 3476 335354 3516
rect 335998 3476 336004 3528
rect 336056 3516 336062 3528
rect 337470 3516 337476 3528
rect 336056 3488 337476 3516
rect 336056 3476 336062 3488
rect 337470 3476 337476 3488
rect 337528 3476 337534 3528
rect 338758 3476 338764 3528
rect 338816 3516 338822 3528
rect 343358 3516 343364 3528
rect 338816 3488 343364 3516
rect 338816 3476 338822 3488
rect 343358 3476 343364 3488
rect 343416 3476 343422 3528
rect 347682 3476 347688 3528
rect 347740 3516 347746 3528
rect 354030 3516 354036 3528
rect 347740 3488 354036 3516
rect 347740 3476 347746 3488
rect 354030 3476 354036 3488
rect 354088 3476 354094 3528
rect 355962 3476 355968 3528
rect 356020 3516 356026 3528
rect 363506 3516 363512 3528
rect 356020 3488 363512 3516
rect 356020 3476 356026 3488
rect 363506 3476 363512 3488
rect 363564 3476 363570 3528
rect 364242 3476 364248 3528
rect 364300 3516 364306 3528
rect 374086 3516 374092 3528
rect 364300 3488 374092 3516
rect 364300 3476 364306 3488
rect 374086 3476 374092 3488
rect 374144 3476 374150 3528
rect 376662 3476 376668 3528
rect 376720 3516 376726 3528
rect 388254 3516 388260 3528
rect 376720 3488 388260 3516
rect 376720 3476 376726 3488
rect 388254 3476 388260 3488
rect 388312 3476 388318 3528
rect 391842 3476 391848 3528
rect 391900 3516 391906 3528
rect 406010 3516 406016 3528
rect 391900 3488 406016 3516
rect 391900 3476 391906 3488
rect 406010 3476 406016 3488
rect 406068 3476 406074 3528
rect 407022 3476 407028 3528
rect 407080 3516 407086 3528
rect 423766 3516 423772 3528
rect 407080 3488 423772 3516
rect 407080 3476 407086 3488
rect 423766 3476 423772 3488
rect 423824 3476 423830 3528
rect 426342 3476 426348 3528
rect 426400 3516 426406 3528
rect 446214 3516 446220 3528
rect 426400 3488 446220 3516
rect 426400 3476 426406 3488
rect 446214 3476 446220 3488
rect 446272 3476 446278 3528
rect 449710 3476 449716 3528
rect 449768 3516 449774 3528
rect 473446 3516 473452 3528
rect 449768 3488 473452 3516
rect 449768 3476 449774 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 476022 3476 476028 3528
rect 476080 3516 476086 3528
rect 504174 3516 504180 3528
rect 476080 3488 504180 3516
rect 476080 3476 476086 3488
rect 504174 3476 504180 3488
rect 504232 3476 504238 3528
rect 506382 3476 506388 3528
rect 506440 3516 506446 3528
rect 538398 3516 538404 3528
rect 506440 3488 538404 3516
rect 506440 3476 506446 3488
rect 538398 3476 538404 3488
rect 538456 3476 538462 3528
rect 539502 3476 539508 3528
rect 539560 3516 539566 3528
rect 577406 3516 577412 3528
rect 539560 3488 577412 3516
rect 539560 3476 539566 3488
rect 577406 3476 577412 3488
rect 577464 3476 577470 3528
rect 128228 3420 132494 3448
rect 128228 3408 128234 3420
rect 134150 3408 134156 3460
rect 134208 3448 134214 3460
rect 135162 3448 135168 3460
rect 134208 3420 135168 3448
rect 134208 3408 134214 3420
rect 135162 3408 135168 3420
rect 135220 3408 135226 3460
rect 138842 3408 138848 3460
rect 138900 3448 138906 3460
rect 139302 3448 139308 3460
rect 138900 3420 139308 3448
rect 138900 3408 138906 3420
rect 139302 3408 139308 3420
rect 139360 3408 139366 3460
rect 141234 3408 141240 3460
rect 141292 3448 141298 3460
rect 142062 3448 142068 3460
rect 141292 3420 142068 3448
rect 141292 3408 141298 3420
rect 142062 3408 142068 3420
rect 142120 3408 142126 3460
rect 161290 3408 161296 3460
rect 161348 3448 161354 3460
rect 180058 3448 180064 3460
rect 161348 3420 180064 3448
rect 161348 3408 161354 3420
rect 180058 3408 180064 3420
rect 180116 3408 180122 3460
rect 189718 3408 189724 3460
rect 189776 3448 189782 3460
rect 190362 3448 190368 3460
rect 189776 3420 190368 3448
rect 189776 3408 189782 3420
rect 190362 3408 190368 3420
rect 190420 3408 190426 3460
rect 265342 3408 265348 3460
rect 265400 3448 265406 3460
rect 266998 3448 267004 3460
rect 265400 3420 267004 3448
rect 265400 3408 265406 3420
rect 266998 3408 267004 3420
rect 267056 3408 267062 3460
rect 272426 3408 272432 3460
rect 272484 3448 272490 3460
rect 273898 3448 273904 3460
rect 272484 3420 273904 3448
rect 272484 3408 272490 3420
rect 273898 3408 273904 3420
rect 273956 3408 273962 3460
rect 321462 3408 321468 3460
rect 321520 3448 321526 3460
rect 323302 3448 323308 3460
rect 321520 3420 323308 3448
rect 321520 3408 321526 3420
rect 323302 3408 323308 3420
rect 323360 3408 323366 3460
rect 325602 3408 325608 3460
rect 325660 3448 325666 3460
rect 329190 3448 329196 3460
rect 325660 3420 329196 3448
rect 325660 3408 325666 3420
rect 329190 3408 329196 3420
rect 329248 3408 329254 3460
rect 331122 3408 331128 3460
rect 331180 3448 331186 3460
rect 335078 3448 335084 3460
rect 331180 3420 335084 3448
rect 331180 3408 331186 3420
rect 335078 3408 335084 3420
rect 335136 3408 335142 3460
rect 335326 3448 335354 3476
rect 339862 3448 339868 3460
rect 335326 3420 339868 3448
rect 339862 3408 339868 3420
rect 339920 3408 339926 3460
rect 342070 3408 342076 3460
rect 342128 3448 342134 3460
rect 348050 3448 348056 3460
rect 342128 3420 348056 3448
rect 342128 3408 342134 3420
rect 348050 3408 348056 3420
rect 348108 3408 348114 3460
rect 361390 3408 361396 3460
rect 361448 3448 361454 3460
rect 370590 3448 370596 3460
rect 361448 3420 370596 3448
rect 361448 3408 361454 3420
rect 370590 3408 370596 3420
rect 370648 3408 370654 3460
rect 372430 3408 372436 3460
rect 372488 3448 372494 3460
rect 383562 3448 383568 3460
rect 372488 3420 383568 3448
rect 372488 3408 372494 3420
rect 383562 3408 383568 3420
rect 383620 3408 383626 3460
rect 383654 3408 383660 3460
rect 383712 3448 383718 3460
rect 396534 3448 396540 3460
rect 383712 3420 396540 3448
rect 383712 3408 383718 3420
rect 396534 3408 396540 3420
rect 396592 3408 396598 3460
rect 398742 3408 398748 3460
rect 398800 3448 398806 3460
rect 414290 3448 414296 3460
rect 398800 3420 414296 3448
rect 398800 3408 398806 3420
rect 414290 3408 414296 3420
rect 414348 3408 414354 3460
rect 417970 3408 417976 3460
rect 418028 3448 418034 3460
rect 436738 3448 436744 3460
rect 418028 3420 436744 3448
rect 418028 3408 418034 3420
rect 436738 3408 436744 3420
rect 436796 3408 436802 3460
rect 445570 3408 445576 3460
rect 445628 3448 445634 3460
rect 468662 3448 468668 3460
rect 445628 3420 468668 3448
rect 445628 3408 445634 3420
rect 468662 3408 468668 3420
rect 468720 3408 468726 3460
rect 469122 3408 469128 3460
rect 469180 3448 469186 3460
rect 495894 3448 495900 3460
rect 469180 3420 495900 3448
rect 469180 3408 469186 3420
rect 495894 3408 495900 3420
rect 495952 3408 495958 3460
rect 499482 3408 499488 3460
rect 499540 3448 499546 3460
rect 530489 3451 530547 3457
rect 530489 3448 530501 3451
rect 499540 3420 530501 3448
rect 499540 3408 499546 3420
rect 530489 3417 530501 3420
rect 530535 3417 530547 3451
rect 530489 3411 530547 3417
rect 530578 3408 530584 3460
rect 530636 3448 530642 3460
rect 536098 3448 536104 3460
rect 530636 3420 536104 3448
rect 530636 3408 530642 3420
rect 536098 3408 536104 3420
rect 536156 3408 536162 3460
rect 548429 3451 548487 3457
rect 548429 3417 548441 3451
rect 548475 3448 548487 3451
rect 552477 3451 552535 3457
rect 552477 3448 552489 3451
rect 548475 3420 552489 3448
rect 548475 3417 548487 3420
rect 548429 3411 548487 3417
rect 552477 3417 552489 3420
rect 552523 3417 552535 3451
rect 552477 3411 552535 3417
rect 552569 3451 552627 3457
rect 552569 3417 552581 3451
rect 552615 3448 552627 3451
rect 582190 3448 582196 3460
rect 552615 3420 582196 3448
rect 552615 3417 552627 3420
rect 552569 3411 552627 3417
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 137278 3380 137284 3392
rect 122806 3352 137284 3380
rect 137278 3340 137284 3352
rect 137336 3340 137342 3392
rect 329650 3340 329656 3392
rect 329708 3380 329714 3392
rect 333882 3380 333888 3392
rect 329708 3352 333888 3380
rect 329708 3340 329714 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 375190 3340 375196 3392
rect 375248 3380 375254 3392
rect 385954 3380 385960 3392
rect 375248 3352 385960 3380
rect 375248 3340 375254 3352
rect 385954 3340 385960 3352
rect 386012 3340 386018 3392
rect 387702 3340 387708 3392
rect 387760 3380 387766 3392
rect 400122 3380 400128 3392
rect 387760 3352 400128 3380
rect 387760 3340 387766 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 401502 3340 401508 3392
rect 401560 3380 401566 3392
rect 416682 3380 416688 3392
rect 401560 3352 416688 3380
rect 401560 3340 401566 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423582 3340 423588 3392
rect 423640 3380 423646 3392
rect 442626 3380 442632 3392
rect 423640 3352 442632 3380
rect 423640 3340 423646 3352
rect 442626 3340 442632 3352
rect 442684 3340 442690 3392
rect 455322 3340 455328 3392
rect 455380 3380 455386 3392
rect 458361 3383 458419 3389
rect 455380 3352 458312 3380
rect 455380 3340 455386 3352
rect 57238 3272 57244 3324
rect 57296 3312 57302 3324
rect 64230 3312 64236 3324
rect 57296 3284 64236 3312
rect 57296 3272 57302 3284
rect 64230 3272 64236 3284
rect 64288 3272 64294 3324
rect 122282 3272 122288 3324
rect 122340 3312 122346 3324
rect 122742 3312 122748 3324
rect 122340 3284 122748 3312
rect 122340 3272 122346 3284
rect 122742 3272 122748 3284
rect 122800 3272 122806 3324
rect 131758 3272 131764 3324
rect 131816 3312 131822 3324
rect 132402 3312 132408 3324
rect 131816 3284 132408 3312
rect 131816 3272 131822 3284
rect 132402 3272 132408 3284
rect 132460 3272 132466 3324
rect 196802 3272 196808 3324
rect 196860 3312 196866 3324
rect 197262 3312 197268 3324
rect 196860 3284 197268 3312
rect 196860 3272 196866 3284
rect 197262 3272 197268 3284
rect 197320 3272 197326 3324
rect 221550 3272 221556 3324
rect 221608 3312 221614 3324
rect 222102 3312 222108 3324
rect 221608 3284 222108 3312
rect 221608 3272 221614 3284
rect 222102 3272 222108 3284
rect 222160 3272 222166 3324
rect 271230 3272 271236 3324
rect 271288 3312 271294 3324
rect 271782 3312 271788 3324
rect 271288 3284 271788 3312
rect 271288 3272 271294 3284
rect 271782 3272 271788 3284
rect 271840 3272 271846 3324
rect 276014 3272 276020 3324
rect 276072 3312 276078 3324
rect 277302 3312 277308 3324
rect 276072 3284 277308 3312
rect 276072 3272 276078 3284
rect 277302 3272 277308 3284
rect 277360 3272 277366 3324
rect 279510 3272 279516 3324
rect 279568 3312 279574 3324
rect 280062 3312 280068 3324
rect 279568 3284 280068 3312
rect 279568 3272 279574 3284
rect 280062 3272 280068 3284
rect 280120 3272 280126 3324
rect 304994 3272 305000 3324
rect 305052 3312 305058 3324
rect 305546 3312 305552 3324
rect 305052 3284 305552 3312
rect 305052 3272 305058 3284
rect 305546 3272 305552 3284
rect 305604 3272 305610 3324
rect 325510 3272 325516 3324
rect 325568 3312 325574 3324
rect 327994 3312 328000 3324
rect 325568 3284 328000 3312
rect 325568 3272 325574 3284
rect 327994 3272 328000 3284
rect 328052 3272 328058 3324
rect 338850 3272 338856 3324
rect 338908 3312 338914 3324
rect 342162 3312 342168 3324
rect 338908 3284 342168 3312
rect 338908 3272 338914 3284
rect 342162 3272 342168 3284
rect 342220 3272 342226 3324
rect 380710 3272 380716 3324
rect 380768 3312 380774 3324
rect 391842 3312 391848 3324
rect 380768 3284 391848 3312
rect 380768 3272 380774 3284
rect 391842 3272 391848 3284
rect 391900 3272 391906 3324
rect 395890 3272 395896 3324
rect 395948 3312 395954 3324
rect 409598 3312 409604 3324
rect 395948 3284 409604 3312
rect 395948 3272 395954 3284
rect 409598 3272 409604 3284
rect 409656 3272 409662 3324
rect 412542 3272 412548 3324
rect 412600 3312 412606 3324
rect 429654 3312 429660 3324
rect 412600 3284 429660 3312
rect 412600 3272 412606 3284
rect 429654 3272 429660 3284
rect 429712 3272 429718 3324
rect 434622 3272 434628 3324
rect 434680 3312 434686 3324
rect 454494 3312 454500 3324
rect 434680 3284 454500 3312
rect 434680 3272 434686 3284
rect 454494 3272 454500 3284
rect 454552 3272 454558 3324
rect 457990 3272 457996 3324
rect 458048 3312 458054 3324
rect 458284 3312 458312 3352
rect 458361 3349 458373 3383
rect 458407 3380 458419 3383
rect 478138 3380 478144 3392
rect 458407 3352 478144 3380
rect 458407 3349 458419 3352
rect 458361 3343 458419 3349
rect 478138 3340 478144 3352
rect 478196 3340 478202 3392
rect 478782 3340 478788 3392
rect 478840 3380 478846 3392
rect 506474 3380 506480 3392
rect 478840 3352 506480 3380
rect 478840 3340 478846 3352
rect 506474 3340 506480 3352
rect 506532 3340 506538 3392
rect 511902 3340 511908 3392
rect 511960 3380 511966 3392
rect 545482 3380 545488 3392
rect 511960 3352 545488 3380
rect 511960 3340 511966 3352
rect 545482 3340 545488 3352
rect 545540 3340 545546 3392
rect 548518 3340 548524 3392
rect 548576 3380 548582 3392
rect 583386 3380 583392 3392
rect 548576 3352 583392 3380
rect 548576 3340 548582 3352
rect 583386 3340 583392 3352
rect 583444 3340 583450 3392
rect 479334 3312 479340 3324
rect 458048 3284 458220 3312
rect 458284 3284 479340 3312
rect 458048 3272 458054 3284
rect 132954 3204 132960 3256
rect 133012 3244 133018 3256
rect 133782 3244 133788 3256
rect 133012 3216 133788 3244
rect 133012 3204 133018 3216
rect 133782 3204 133788 3216
rect 133840 3204 133846 3256
rect 183738 3204 183744 3256
rect 183796 3244 183802 3256
rect 184842 3244 184848 3256
rect 183796 3216 184848 3244
rect 183796 3204 183802 3216
rect 184842 3204 184848 3216
rect 184900 3204 184906 3256
rect 200298 3204 200304 3256
rect 200356 3244 200362 3256
rect 201402 3244 201408 3256
rect 200356 3216 201408 3244
rect 200356 3204 200362 3216
rect 201402 3204 201408 3216
rect 201460 3204 201466 3256
rect 225138 3204 225144 3256
rect 225196 3244 225202 3256
rect 226242 3244 226248 3256
rect 225196 3216 226248 3244
rect 225196 3204 225202 3216
rect 226242 3204 226248 3216
rect 226300 3204 226306 3256
rect 309134 3204 309140 3256
rect 309192 3244 309198 3256
rect 310238 3244 310244 3256
rect 309192 3216 310244 3244
rect 309192 3204 309198 3216
rect 310238 3204 310244 3216
rect 310296 3204 310302 3256
rect 322842 3204 322848 3256
rect 322900 3244 322906 3256
rect 325602 3244 325608 3256
rect 322900 3216 325608 3244
rect 322900 3204 322906 3216
rect 325602 3204 325608 3216
rect 325660 3204 325666 3256
rect 336642 3204 336648 3256
rect 336700 3244 336706 3256
rect 340966 3244 340972 3256
rect 336700 3216 340972 3244
rect 336700 3204 336706 3216
rect 340966 3204 340972 3216
rect 341024 3204 341030 3256
rect 402882 3204 402888 3256
rect 402940 3244 402946 3256
rect 417878 3244 417884 3256
rect 402940 3216 417884 3244
rect 402940 3204 402946 3216
rect 417878 3204 417884 3216
rect 417936 3204 417942 3256
rect 418062 3204 418068 3256
rect 418120 3244 418126 3256
rect 435542 3244 435548 3256
rect 418120 3216 435548 3244
rect 418120 3204 418126 3216
rect 435542 3204 435548 3216
rect 435600 3204 435606 3256
rect 437382 3204 437388 3256
rect 437440 3244 437446 3256
rect 458082 3244 458088 3256
rect 437440 3216 458088 3244
rect 437440 3204 437446 3216
rect 458082 3204 458088 3216
rect 458140 3204 458146 3256
rect 458192 3244 458220 3284
rect 479334 3272 479340 3284
rect 479392 3272 479398 3324
rect 481542 3272 481548 3324
rect 481600 3312 481606 3324
rect 510062 3312 510068 3324
rect 481600 3284 510068 3312
rect 481600 3272 481606 3284
rect 510062 3272 510068 3284
rect 510120 3272 510126 3324
rect 514662 3272 514668 3324
rect 514720 3312 514726 3324
rect 549070 3312 549076 3324
rect 514720 3284 549076 3312
rect 514720 3272 514726 3284
rect 549070 3272 549076 3284
rect 549128 3272 549134 3324
rect 549162 3272 549168 3324
rect 549220 3312 549226 3324
rect 580994 3312 581000 3324
rect 549220 3284 581000 3312
rect 549220 3272 549226 3284
rect 580994 3272 581000 3284
rect 581052 3272 581058 3324
rect 482830 3244 482836 3256
rect 458192 3216 482836 3244
rect 482830 3204 482836 3216
rect 482888 3204 482894 3256
rect 488442 3204 488448 3256
rect 488500 3244 488506 3256
rect 517146 3244 517152 3256
rect 488500 3216 517152 3244
rect 488500 3204 488506 3216
rect 517146 3204 517152 3216
rect 517204 3204 517210 3256
rect 522942 3204 522948 3256
rect 523000 3244 523006 3256
rect 557350 3244 557356 3256
rect 523000 3216 557356 3244
rect 523000 3204 523006 3216
rect 557350 3204 557356 3216
rect 557408 3204 557414 3256
rect 241698 3136 241704 3188
rect 241756 3176 241762 3188
rect 242802 3176 242808 3188
rect 241756 3148 242808 3176
rect 241756 3136 241762 3148
rect 242802 3136 242808 3148
rect 242860 3136 242866 3188
rect 283098 3136 283104 3188
rect 283156 3176 283162 3188
rect 285766 3176 285772 3188
rect 283156 3148 285772 3176
rect 283156 3136 283162 3148
rect 285766 3136 285772 3148
rect 285824 3136 285830 3188
rect 326982 3136 326988 3188
rect 327040 3176 327046 3188
rect 330386 3176 330392 3188
rect 327040 3148 330392 3176
rect 327040 3136 327046 3148
rect 330386 3136 330392 3148
rect 330444 3136 330450 3188
rect 390462 3136 390468 3188
rect 390520 3176 390526 3188
rect 403618 3176 403624 3188
rect 390520 3148 403624 3176
rect 390520 3136 390526 3148
rect 403618 3136 403624 3148
rect 403676 3136 403682 3188
rect 408310 3136 408316 3188
rect 408368 3176 408374 3188
rect 408368 3148 412634 3176
rect 408368 3136 408374 3148
rect 246390 3068 246396 3120
rect 246448 3108 246454 3120
rect 246942 3108 246948 3120
rect 246448 3080 246948 3108
rect 246448 3068 246454 3080
rect 246942 3068 246948 3080
rect 247000 3068 247006 3120
rect 297266 3068 297272 3120
rect 297324 3108 297330 3120
rect 298186 3108 298192 3120
rect 297324 3080 298192 3108
rect 297324 3068 297330 3080
rect 298186 3068 298192 3080
rect 298244 3068 298250 3120
rect 394602 3068 394608 3120
rect 394660 3108 394666 3120
rect 408402 3108 408408 3120
rect 394660 3080 408408 3108
rect 394660 3068 394666 3080
rect 408402 3068 408408 3080
rect 408460 3068 408466 3120
rect 412606 3108 412634 3148
rect 420822 3136 420828 3188
rect 420880 3176 420886 3188
rect 439130 3176 439136 3188
rect 420880 3148 439136 3176
rect 420880 3136 420886 3148
rect 439130 3136 439136 3148
rect 439188 3136 439194 3188
rect 453850 3136 453856 3188
rect 453908 3176 453914 3188
rect 476942 3176 476948 3188
rect 453908 3148 476948 3176
rect 453908 3136 453914 3148
rect 476942 3136 476948 3148
rect 477000 3136 477006 3188
rect 482922 3136 482928 3188
rect 482980 3176 482986 3188
rect 511258 3176 511264 3188
rect 482980 3148 511264 3176
rect 482980 3136 482986 3148
rect 511258 3136 511264 3148
rect 511316 3136 511322 3188
rect 516042 3136 516048 3188
rect 516100 3176 516106 3188
rect 550266 3176 550272 3188
rect 516100 3148 550272 3176
rect 516100 3136 516106 3148
rect 550266 3136 550272 3148
rect 550324 3136 550330 3188
rect 552477 3179 552535 3185
rect 552477 3145 552489 3179
rect 552523 3176 552535 3179
rect 556154 3176 556160 3188
rect 552523 3148 556160 3176
rect 552523 3145 552535 3148
rect 552477 3139 552535 3145
rect 556154 3136 556160 3148
rect 556212 3136 556218 3188
rect 424962 3108 424968 3120
rect 412606 3080 424968 3108
rect 424962 3068 424968 3080
rect 425020 3068 425026 3120
rect 430482 3068 430488 3120
rect 430540 3108 430546 3120
rect 449802 3108 449808 3120
rect 430540 3080 449808 3108
rect 430540 3068 430546 3080
rect 449802 3068 449808 3080
rect 449860 3068 449866 3120
rect 451182 3068 451188 3120
rect 451240 3108 451246 3120
rect 474550 3108 474556 3120
rect 451240 3080 474556 3108
rect 451240 3068 451246 3080
rect 474550 3068 474556 3080
rect 474608 3068 474614 3120
rect 480162 3068 480168 3120
rect 480220 3108 480226 3120
rect 507670 3108 507676 3120
rect 480220 3080 507676 3108
rect 480220 3068 480226 3080
rect 507670 3068 507676 3080
rect 507728 3068 507734 3120
rect 513282 3068 513288 3120
rect 513340 3108 513346 3120
rect 546678 3108 546684 3120
rect 513340 3080 546684 3108
rect 513340 3068 513346 3080
rect 546678 3068 546684 3080
rect 546736 3068 546742 3120
rect 547138 3068 547144 3120
rect 547196 3108 547202 3120
rect 578602 3108 578608 3120
rect 547196 3080 578608 3108
rect 547196 3068 547202 3080
rect 578602 3068 578608 3080
rect 578660 3068 578666 3120
rect 135254 3000 135260 3052
rect 135312 3040 135318 3052
rect 136542 3040 136548 3052
rect 135312 3012 136548 3040
rect 135312 3000 135318 3012
rect 136542 3000 136548 3012
rect 136600 3000 136606 3052
rect 140038 3000 140044 3052
rect 140096 3040 140102 3052
rect 140682 3040 140688 3052
rect 140096 3012 140688 3040
rect 140096 3000 140102 3012
rect 140682 3000 140688 3012
rect 140740 3000 140746 3052
rect 164878 3000 164884 3052
rect 164936 3040 164942 3052
rect 165522 3040 165528 3052
rect 164936 3012 165528 3040
rect 164936 3000 164942 3012
rect 165522 3000 165528 3012
rect 165580 3000 165586 3052
rect 201494 3000 201500 3052
rect 201552 3040 201558 3052
rect 202598 3040 202604 3052
rect 201552 3012 202604 3040
rect 201552 3000 201558 3012
rect 202598 3000 202604 3012
rect 202656 3000 202662 3052
rect 208578 3000 208584 3052
rect 208636 3040 208642 3052
rect 209682 3040 209688 3052
rect 208636 3012 209688 3040
rect 208636 3000 208642 3012
rect 209682 3000 209688 3012
rect 209740 3000 209746 3052
rect 248782 3000 248788 3052
rect 248840 3040 248846 3052
rect 249702 3040 249708 3052
rect 248840 3012 249708 3040
rect 248840 3000 248846 3012
rect 249702 3000 249708 3012
rect 249760 3000 249766 3052
rect 318610 3000 318616 3052
rect 318668 3040 318674 3052
rect 320910 3040 320916 3052
rect 318668 3012 320916 3040
rect 318668 3000 318674 3012
rect 320910 3000 320916 3012
rect 320968 3000 320974 3052
rect 346302 3000 346308 3052
rect 346360 3040 346366 3052
rect 352834 3040 352840 3052
rect 346360 3012 352840 3040
rect 346360 3000 346366 3012
rect 352834 3000 352840 3012
rect 352892 3000 352898 3052
rect 416590 3000 416596 3052
rect 416648 3040 416654 3052
rect 434438 3040 434444 3052
rect 416648 3012 434444 3040
rect 416648 3000 416654 3012
rect 434438 3000 434444 3012
rect 434496 3000 434502 3052
rect 445662 3000 445668 3052
rect 445720 3040 445726 3052
rect 467466 3040 467472 3052
rect 445720 3012 467472 3040
rect 445720 3000 445726 3012
rect 467466 3000 467472 3012
rect 467524 3000 467530 3052
rect 473262 3000 473268 3052
rect 473320 3040 473326 3052
rect 500586 3040 500592 3052
rect 473320 3012 500592 3040
rect 473320 3000 473326 3012
rect 500586 3000 500592 3012
rect 500644 3000 500650 3052
rect 509142 3000 509148 3052
rect 509200 3040 509206 3052
rect 541986 3040 541992 3052
rect 509200 3012 541992 3040
rect 509200 3000 509206 3012
rect 541986 3000 541992 3012
rect 542044 3000 542050 3052
rect 542262 3000 542268 3052
rect 542320 3040 542326 3052
rect 552569 3043 552627 3049
rect 552569 3040 552581 3043
rect 542320 3012 552581 3040
rect 542320 3000 542326 3012
rect 552569 3009 552581 3012
rect 552615 3009 552627 3043
rect 552569 3003 552627 3009
rect 552661 3043 552719 3049
rect 552661 3009 552673 3043
rect 552707 3040 552719 3043
rect 571518 3040 571524 3052
rect 552707 3012 571524 3040
rect 552707 3009 552719 3012
rect 552661 3003 552719 3009
rect 571518 3000 571524 3012
rect 571576 3000 571582 3052
rect 320818 2932 320824 2984
rect 320876 2972 320882 2984
rect 322106 2972 322112 2984
rect 320876 2944 322112 2972
rect 320876 2932 320882 2944
rect 322106 2932 322112 2944
rect 322164 2932 322170 2984
rect 349062 2932 349068 2984
rect 349120 2972 349126 2984
rect 356330 2972 356336 2984
rect 349120 2944 356336 2972
rect 349120 2932 349126 2944
rect 356330 2932 356336 2944
rect 356388 2932 356394 2984
rect 413922 2932 413928 2984
rect 413980 2972 413986 2984
rect 430850 2972 430856 2984
rect 413980 2944 430856 2972
rect 413980 2932 413986 2944
rect 430850 2932 430856 2944
rect 430908 2932 430914 2984
rect 440142 2932 440148 2984
rect 440200 2972 440206 2984
rect 461578 2972 461584 2984
rect 440200 2944 461584 2972
rect 440200 2932 440206 2944
rect 461578 2932 461584 2944
rect 461636 2932 461642 2984
rect 466362 2932 466368 2984
rect 466420 2972 466426 2984
rect 492306 2972 492312 2984
rect 466420 2944 492312 2972
rect 466420 2932 466426 2944
rect 492306 2932 492312 2944
rect 492364 2932 492370 2984
rect 497458 2932 497464 2984
rect 497516 2972 497522 2984
rect 518342 2972 518348 2984
rect 497516 2944 518348 2972
rect 497516 2932 497522 2944
rect 518342 2932 518348 2944
rect 518400 2932 518406 2984
rect 530489 2975 530547 2981
rect 530489 2941 530501 2975
rect 530535 2972 530547 2975
rect 531314 2972 531320 2984
rect 530535 2944 531320 2972
rect 530535 2941 530547 2944
rect 530489 2935 530547 2941
rect 531314 2932 531320 2944
rect 531372 2932 531378 2984
rect 540238 2932 540244 2984
rect 540296 2972 540302 2984
rect 564434 2972 564440 2984
rect 540296 2944 564440 2972
rect 540296 2932 540302 2944
rect 564434 2932 564440 2944
rect 564492 2932 564498 2984
rect 65518 2864 65524 2916
rect 65576 2904 65582 2916
rect 66162 2904 66168 2916
rect 65576 2876 66168 2904
rect 65576 2864 65582 2876
rect 66162 2864 66168 2876
rect 66220 2864 66226 2916
rect 409782 2864 409788 2916
rect 409840 2904 409846 2916
rect 426158 2904 426164 2916
rect 409840 2876 426164 2904
rect 409840 2864 409846 2876
rect 426158 2864 426164 2876
rect 426216 2864 426222 2916
rect 444282 2864 444288 2916
rect 444340 2904 444346 2916
rect 466270 2904 466276 2916
rect 444340 2876 466276 2904
rect 444340 2864 444346 2876
rect 466270 2864 466276 2876
rect 466328 2864 466334 2916
rect 545758 2864 545764 2916
rect 545816 2904 545822 2916
rect 552661 2907 552719 2913
rect 552661 2904 552673 2907
rect 545816 2876 552673 2904
rect 545816 2864 545822 2876
rect 552661 2873 552673 2876
rect 552707 2873 552719 2907
rect 568022 2904 568028 2916
rect 552661 2867 552719 2873
rect 557506 2876 568028 2904
rect 294874 2796 294880 2848
rect 294932 2836 294938 2848
rect 295426 2836 295432 2848
rect 294932 2808 295432 2836
rect 294932 2796 294938 2808
rect 295426 2796 295432 2808
rect 295484 2796 295490 2848
rect 454678 2796 454684 2848
rect 454736 2836 454742 2848
rect 475746 2836 475752 2848
rect 454736 2808 475752 2836
rect 454736 2796 454742 2808
rect 475746 2796 475752 2808
rect 475804 2796 475810 2848
rect 544470 2796 544476 2848
rect 544528 2836 544534 2848
rect 557506 2836 557534 2876
rect 568022 2864 568028 2876
rect 568080 2864 568086 2916
rect 544528 2808 557534 2836
rect 544528 2796 544534 2808
<< via1 >>
rect 154120 700952 154172 701004
rect 329840 700952 329892 701004
rect 137836 700884 137888 700936
rect 325700 700884 325752 700936
rect 336004 700884 336056 700936
rect 364984 700884 365036 700936
rect 260748 700816 260800 700868
rect 462320 700816 462372 700868
rect 264888 700748 264940 700800
rect 478512 700748 478564 700800
rect 89168 700680 89220 700732
rect 343640 700680 343692 700732
rect 72976 700612 73028 700664
rect 338120 700612 338172 700664
rect 340144 700612 340196 700664
rect 494796 700612 494848 700664
rect 246948 700544 247000 700596
rect 527180 700544 527232 700596
rect 252468 700476 252520 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 347780 700408 347832 700460
rect 24308 700340 24360 700392
rect 356060 700340 356112 700392
rect 8116 700272 8168 700324
rect 351920 700272 351972 700324
rect 543004 700272 543056 700324
rect 559656 700272 559708 700324
rect 278688 700204 278740 700256
rect 413652 700204 413704 700256
rect 274548 700136 274600 700188
rect 397460 700136 397512 700188
rect 202788 700068 202840 700120
rect 311900 700068 311952 700120
rect 218980 700000 219032 700052
rect 316040 700000 316092 700052
rect 291108 699932 291160 699984
rect 348792 699932 348844 699984
rect 286968 699864 287020 699916
rect 332508 699864 332560 699916
rect 267648 699796 267700 699848
rect 299572 699796 299624 699848
rect 283840 699728 283892 699780
rect 303620 699728 303672 699780
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 173164 699660 173216 699712
rect 235172 699660 235224 699712
rect 240784 699660 240836 699712
rect 296628 698912 296680 698964
rect 300124 698912 300176 698964
rect 234528 696940 234580 696992
rect 580172 696940 580224 696992
rect 238668 683204 238720 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 360200 683136 360252 683188
rect 229836 670760 229888 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 369860 670692 369912 670744
rect 282092 660288 282144 660340
rect 336004 660288 336056 660340
rect 240784 659268 240836 659320
rect 308496 659268 308548 659320
rect 255780 659200 255832 659252
rect 340144 659200 340196 659252
rect 173164 659132 173216 659184
rect 321652 659132 321704 659184
rect 268936 659064 268988 659116
rect 429200 659064 429252 659116
rect 106188 658996 106240 659048
rect 334808 658996 334860 659048
rect 242532 658928 242584 658980
rect 543004 658928 543056 658980
rect 29644 658316 29696 658368
rect 541348 658316 541400 658368
rect 53656 658248 53708 658300
rect 566464 658248 566516 658300
rect 211804 658180 211856 658232
rect 565176 658180 565228 658232
rect 194232 658112 194284 658164
rect 548616 658112 548668 658164
rect 3424 658044 3476 658096
rect 365628 658044 365680 658096
rect 42248 657976 42300 658028
rect 409512 657976 409564 658028
rect 132776 657908 132828 657960
rect 184848 657908 184900 657960
rect 185492 657908 185544 657960
rect 556896 657908 556948 657960
rect 167920 657840 167972 657892
rect 551376 657840 551428 657892
rect 181076 657772 181128 657824
rect 576216 657772 576268 657824
rect 25596 657704 25648 657756
rect 435916 657704 435968 657756
rect 163504 657636 163556 657688
rect 573456 657636 573508 657688
rect 154672 657568 154724 657620
rect 574836 657568 574888 657620
rect 137100 657500 137152 657552
rect 566556 657500 566608 657552
rect 39304 657432 39356 657484
rect 471060 657432 471112 657484
rect 36544 657364 36596 657416
rect 475384 657364 475436 657416
rect 11704 657296 11756 657348
rect 462228 657296 462280 657348
rect 110788 657228 110840 657280
rect 562416 657228 562468 657280
rect 42064 657160 42116 657212
rect 501788 657160 501840 657212
rect 88800 657092 88852 657144
rect 548524 657092 548576 657144
rect 15844 657024 15896 657076
rect 484216 657024 484268 657076
rect 75644 656956 75696 657008
rect 545764 656956 545816 657008
rect 84384 656888 84436 656940
rect 558184 656888 558236 656940
rect 216220 656820 216272 656872
rect 548708 656820 548760 656872
rect 203064 656752 203116 656804
rect 547236 656752 547288 656804
rect 189816 656684 189868 656736
rect 545856 656684 545908 656736
rect 11888 656616 11940 656668
rect 374368 656616 374420 656668
rect 176660 656548 176712 656600
rect 544476 656548 544528 656600
rect 14556 656480 14608 656532
rect 387524 656480 387576 656532
rect 15936 656412 15988 656464
rect 400772 656412 400824 656464
rect 17316 656344 17368 656396
rect 413928 656344 413980 656396
rect 159088 656276 159140 656328
rect 555516 656276 555568 656328
rect 18696 656208 18748 656260
rect 427084 656208 427136 656260
rect 172244 656140 172296 656192
rect 580356 656140 580408 656192
rect 21456 656072 21508 656124
rect 440240 656072 440292 656124
rect 22744 656004 22796 656056
rect 453488 656004 453540 656056
rect 25504 655936 25556 655988
rect 466644 655936 466696 655988
rect 123944 655868 123996 655920
rect 565084 655868 565136 655920
rect 29736 655800 29788 655852
rect 492956 655800 493008 655852
rect 97632 655732 97684 655784
rect 561036 655732 561088 655784
rect 7564 655664 7616 655716
rect 479524 655664 479576 655716
rect 32404 655596 32456 655648
rect 505836 655596 505888 655648
rect 71504 655528 71556 655580
rect 556804 655528 556856 655580
rect 184848 655392 184900 655444
rect 580264 655392 580316 655444
rect 225328 655324 225380 655376
rect 558368 655324 558420 655376
rect 102140 655299 102192 655308
rect 102140 655265 102149 655299
rect 102149 655265 102183 655299
rect 102183 655265 102192 655299
rect 102140 655256 102192 655265
rect 106648 655299 106700 655308
rect 106648 655265 106657 655299
rect 106657 655265 106691 655299
rect 106691 655265 106700 655299
rect 106648 655256 106700 655265
rect 115480 655299 115532 655308
rect 115480 655265 115489 655299
rect 115489 655265 115523 655299
rect 115523 655265 115532 655299
rect 115480 655256 115532 655265
rect 119896 655299 119948 655308
rect 119896 655265 119905 655299
rect 119905 655265 119939 655299
rect 119939 655265 119948 655299
rect 119896 655256 119948 655265
rect 128728 655299 128780 655308
rect 128728 655265 128737 655299
rect 128737 655265 128771 655299
rect 128771 655265 128780 655299
rect 128728 655256 128780 655265
rect 141792 655299 141844 655308
rect 141792 655265 141801 655299
rect 141801 655265 141835 655299
rect 141835 655265 141844 655299
rect 141792 655256 141844 655265
rect 146208 655299 146260 655308
rect 146208 655265 146217 655299
rect 146217 655265 146251 655299
rect 146251 655265 146260 655299
rect 146208 655256 146260 655265
rect 198556 655256 198608 655308
rect 554044 655256 554096 655308
rect 40776 655188 40828 655240
rect 404820 655188 404872 655240
rect 7656 655120 7708 655172
rect 382924 655120 382976 655172
rect 42156 655052 42208 655104
rect 418160 655052 418212 655104
rect 10324 654984 10376 655036
rect 396080 654984 396132 655036
rect 22836 654916 22888 654968
rect 422484 654984 422536 655036
rect 431132 655027 431184 655036
rect 431132 654993 431141 655027
rect 431141 654993 431175 655027
rect 431175 654993 431184 655027
rect 431132 654984 431184 654993
rect 444380 654984 444432 655036
rect 448796 655027 448848 655036
rect 448796 654993 448805 655027
rect 448805 654993 448839 655027
rect 448839 654993 448848 655027
rect 448796 654984 448848 654993
rect 457444 655027 457496 655036
rect 457444 654993 457453 655027
rect 457453 654993 457487 655027
rect 457487 654993 457496 655027
rect 457444 654984 457496 654993
rect 488540 655027 488592 655036
rect 488540 654993 488549 655027
rect 488549 654993 488583 655027
rect 488583 654993 488592 655027
rect 488540 654984 488592 654993
rect 36636 654848 36688 654900
rect 558276 654780 558328 654832
rect 11796 654712 11848 654764
rect 26884 654644 26936 654696
rect 569224 654576 569276 654628
rect 544384 654508 544436 654560
rect 14464 654440 14516 654492
rect 573364 654372 573416 654424
rect 578884 654304 578936 654356
rect 571984 654236 572036 654288
rect 576124 654168 576176 654220
rect 3516 654100 3568 654152
rect 561128 644376 561180 644428
rect 580172 644376 580224 644428
rect 3332 633360 3384 633412
rect 11888 633360 11940 633412
rect 558368 632000 558420 632052
rect 580172 632000 580224 632052
rect 3148 619284 3200 619336
rect 7656 619284 7708 619336
rect 548708 618196 548760 618248
rect 580172 618196 580224 618248
rect 3056 607112 3108 607164
rect 36728 607112 36780 607164
rect 555608 591948 555660 592000
rect 580172 591948 580224 592000
rect 3332 580932 3384 580984
rect 14556 580932 14608 580984
rect 565176 578144 565228 578196
rect 579620 578144 579672 578196
rect 3332 567128 3384 567180
rect 10324 567128 10376 567180
rect 547236 564340 547288 564392
rect 580172 564340 580224 564392
rect 3332 554684 3384 554736
rect 39396 554684 39448 554736
rect 548616 538160 548668 538212
rect 580172 538160 580224 538212
rect 3332 528504 3384 528556
rect 15936 528504 15988 528556
rect 554044 525716 554096 525768
rect 579896 525716 579948 525768
rect 3148 516060 3200 516112
rect 42248 516060 42300 516112
rect 545856 511912 545908 511964
rect 580172 511912 580224 511964
rect 2964 502256 3016 502308
rect 40776 502256 40828 502308
rect 576216 485732 576268 485784
rect 580172 485732 580224 485784
rect 3240 476008 3292 476060
rect 17316 476008 17368 476060
rect 556896 471928 556948 471980
rect 579620 471928 579672 471980
rect 3056 463632 3108 463684
rect 22836 463632 22888 463684
rect 544476 458124 544528 458176
rect 580172 458124 580224 458176
rect 3332 449828 3384 449880
rect 42156 449828 42208 449880
rect 551376 431876 551428 431928
rect 579620 431876 579672 431928
rect 3332 423580 3384 423632
rect 18696 423580 18748 423632
rect 2964 411204 3016 411256
rect 25596 411204 25648 411256
rect 573456 405628 573508 405680
rect 579620 405628 579672 405680
rect 3332 398760 3384 398812
rect 11796 398760 11848 398812
rect 574836 379448 574888 379500
rect 580172 379448 580224 379500
rect 3332 372512 3384 372564
rect 21456 372512 21508 372564
rect 555516 365644 555568 365696
rect 580172 365644 580224 365696
rect 3332 358708 3384 358760
rect 26884 358708 26936 358760
rect 569316 353200 569368 353252
rect 580172 353200 580224 353252
rect 3332 346332 3384 346384
rect 36636 346332 36688 346384
rect 569224 325592 569276 325644
rect 579896 325592 579948 325644
rect 3332 320084 3384 320136
rect 22744 320084 22796 320136
rect 558276 313216 558328 313268
rect 580172 313216 580224 313268
rect 3332 306280 3384 306332
rect 11704 306280 11756 306332
rect 566556 299412 566608 299464
rect 579620 299412 579672 299464
rect 3332 293904 3384 293956
rect 14464 293904 14516 293956
rect 573364 273164 573416 273216
rect 579896 273164 579948 273216
rect 2964 267656 3016 267708
rect 25504 267656 25556 267708
rect 3148 255212 3200 255264
rect 36544 255212 36596 255264
rect 565084 245556 565136 245608
rect 580172 245556 580224 245608
rect 3240 241408 3292 241460
rect 39304 241408 39356 241460
rect 544384 233180 544436 233232
rect 579988 233180 580040 233232
rect 3332 214956 3384 215008
rect 7564 214956 7616 215008
rect 562416 206932 562468 206984
rect 579804 206932 579856 206984
rect 576124 193128 576176 193180
rect 580172 193128 580224 193180
rect 3516 188980 3568 189032
rect 15844 188980 15896 189032
rect 571984 179324 572036 179376
rect 580172 179324 580224 179376
rect 561036 166948 561088 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 29736 164160 29788 164212
rect 548524 153144 548576 153196
rect 580172 153144 580224 153196
rect 3516 150356 3568 150408
rect 42064 150356 42116 150408
rect 570604 139340 570656 139392
rect 580172 139340 580224 139392
rect 3516 137912 3568 137964
rect 40684 137912 40736 137964
rect 558184 126896 558236 126948
rect 580172 126896 580224 126948
rect 545764 113092 545816 113144
rect 579804 113092 579856 113144
rect 3148 111732 3200 111784
rect 32404 111732 32456 111784
rect 560944 100648 560996 100700
rect 580172 100648 580224 100700
rect 556804 86912 556856 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 17224 85484 17276 85536
rect 547144 73108 547196 73160
rect 580172 73108 580224 73160
rect 3424 71680 3476 71732
rect 33784 71680 33836 71732
rect 562324 60664 562376 60716
rect 580172 60664 580224 60716
rect 2780 58624 2832 58676
rect 4804 58624 4856 58676
rect 23388 51008 23440 51060
rect 62488 51008 62540 51060
rect 71044 51008 71096 51060
rect 81808 51008 81860 51060
rect 19248 50940 19300 50992
rect 58440 50940 58492 50992
rect 16488 50872 16540 50924
rect 56416 50872 56468 50924
rect 57244 50872 57296 50924
rect 78772 50940 78824 50992
rect 81348 50940 81400 50992
rect 112260 51008 112312 51060
rect 115848 51008 115900 51060
rect 141792 51008 141844 51060
rect 144644 51008 144696 51060
rect 166172 51008 166224 51060
rect 168288 51008 168340 51060
rect 186504 51008 186556 51060
rect 190368 51008 190420 51060
rect 205732 51008 205784 51060
rect 208308 51008 208360 51060
rect 221004 51008 221056 51060
rect 222108 51008 222160 51060
rect 233148 51008 233200 51060
rect 530860 51008 530912 51060
rect 544384 51008 544436 51060
rect 109224 50940 109276 50992
rect 113088 50940 113140 50992
rect 139768 50940 139820 50992
rect 140688 50940 140740 50992
rect 163136 50940 163188 50992
rect 182364 50940 182416 50992
rect 183468 50940 183520 50992
rect 199660 50940 199712 50992
rect 200028 50940 200080 50992
rect 213920 50940 213972 50992
rect 215208 50940 215260 50992
rect 227076 50940 227128 50992
rect 227628 50940 227680 50992
rect 237288 50940 237340 50992
rect 241428 50940 241480 50992
rect 249432 50940 249484 50992
rect 252376 50940 252428 50992
rect 259644 50940 259696 50992
rect 510528 50940 510580 50992
rect 536104 50940 536156 50992
rect 67548 50872 67600 50924
rect 12348 50804 12400 50856
rect 52368 50804 52420 50856
rect 56508 50804 56560 50856
rect 67640 50804 67692 50856
rect 20628 50736 20680 50788
rect 59452 50736 59504 50788
rect 63408 50736 63460 50788
rect 70308 50872 70360 50924
rect 103152 50872 103204 50924
rect 110328 50872 110380 50924
rect 136640 50872 136692 50924
rect 139308 50872 139360 50924
rect 162032 50872 162084 50924
rect 165528 50872 165580 50924
rect 184388 50872 184440 50924
rect 186228 50872 186280 50924
rect 201684 50872 201736 50924
rect 205548 50872 205600 50924
rect 218980 50872 219032 50924
rect 219256 50872 219308 50924
rect 230112 50872 230164 50924
rect 234528 50872 234580 50924
rect 243360 50872 243412 50924
rect 253848 50872 253900 50924
rect 260656 50872 260708 50924
rect 509516 50872 509568 50924
rect 542360 50872 542412 50924
rect 68928 50804 68980 50856
rect 101128 50804 101180 50856
rect 107568 50804 107620 50856
rect 134616 50804 134668 50856
rect 144736 50804 144788 50856
rect 167184 50804 167236 50856
rect 179328 50804 179380 50856
rect 180064 50804 180116 50856
rect 10968 50668 11020 50720
rect 51356 50668 51408 50720
rect 54484 50668 54536 50720
rect 63500 50668 63552 50720
rect 15108 50600 15160 50652
rect 55404 50600 55456 50652
rect 55864 50600 55916 50652
rect 13728 50532 13780 50584
rect 54392 50532 54444 50584
rect 60648 50532 60700 50584
rect 66536 50600 66588 50652
rect 100116 50736 100168 50788
rect 103428 50736 103480 50788
rect 130568 50736 130620 50788
rect 137928 50736 137980 50788
rect 161020 50736 161072 50788
rect 161388 50736 161440 50788
rect 180340 50736 180392 50788
rect 190552 50804 190604 50856
rect 194416 50804 194468 50856
rect 208768 50804 208820 50856
rect 211068 50804 211120 50856
rect 223028 50804 223080 50856
rect 223488 50804 223540 50856
rect 234252 50804 234304 50856
rect 235908 50804 235960 50856
rect 244372 50804 244424 50856
rect 262128 50804 262180 50856
rect 267740 50804 267792 50856
rect 506480 50804 506532 50856
rect 543004 50804 543056 50856
rect 548524 50804 548576 50856
rect 181352 50736 181404 50788
rect 89076 50668 89128 50720
rect 95056 50668 95108 50720
rect 95148 50668 95200 50720
rect 99288 50668 99340 50720
rect 127532 50668 127584 50720
rect 136548 50668 136600 50720
rect 158996 50668 159048 50720
rect 160008 50668 160060 50720
rect 166908 50668 166960 50720
rect 185400 50668 185452 50720
rect 97080 50600 97132 50652
rect 100668 50600 100720 50652
rect 128544 50600 128596 50652
rect 135168 50600 135220 50652
rect 157984 50600 158036 50652
rect 162768 50600 162820 50652
rect 180708 50600 180760 50652
rect 197636 50736 197688 50788
rect 198648 50736 198700 50788
rect 212908 50736 212960 50788
rect 213828 50736 213880 50788
rect 226064 50736 226116 50788
rect 226248 50736 226300 50788
rect 236276 50736 236328 50788
rect 237288 50736 237340 50788
rect 246396 50736 246448 50788
rect 246948 50736 247000 50788
rect 254492 50736 254544 50788
rect 264888 50736 264940 50788
rect 269764 50736 269816 50788
rect 275928 50736 275980 50788
rect 278872 50736 278924 50788
rect 285496 50736 285548 50788
rect 288072 50736 288124 50788
rect 332784 50736 332836 50788
rect 336004 50736 336056 50788
rect 458732 50736 458784 50788
rect 461584 50736 461636 50788
rect 477040 50736 477092 50788
rect 482284 50736 482336 50788
rect 516600 50736 516652 50788
rect 520924 50736 520976 50788
rect 522764 50736 522816 50788
rect 556804 50736 556856 50788
rect 187608 50668 187660 50720
rect 203708 50668 203760 50720
rect 204168 50668 204220 50720
rect 217968 50668 218020 50720
rect 219348 50668 219400 50720
rect 231124 50668 231176 50720
rect 231768 50668 231820 50720
rect 241336 50668 241388 50720
rect 244188 50668 244240 50720
rect 252468 50668 252520 50720
rect 267648 50668 267700 50720
rect 271788 50668 271840 50720
rect 277308 50668 277360 50720
rect 279884 50668 279936 50720
rect 285588 50668 285640 50720
rect 287060 50668 287112 50720
rect 525800 50668 525852 50720
rect 560944 50668 560996 50720
rect 186136 50600 186188 50652
rect 202696 50600 202748 50652
rect 202788 50600 202840 50652
rect 215944 50600 215996 50652
rect 216588 50600 216640 50652
rect 228088 50600 228140 50652
rect 229008 50600 229060 50652
rect 239312 50600 239364 50652
rect 240048 50600 240100 50652
rect 248420 50600 248472 50652
rect 256608 50600 256660 50652
rect 262680 50600 262732 50652
rect 274548 50600 274600 50652
rect 277860 50600 277912 50652
rect 492220 50600 492272 50652
rect 500224 50600 500276 50652
rect 528836 50600 528888 50652
rect 564532 50600 564584 50652
rect 91008 50532 91060 50584
rect 9588 50464 9640 50516
rect 50344 50464 50396 50516
rect 53748 50464 53800 50516
rect 87880 50464 87932 50516
rect 6828 50396 6880 50448
rect 48320 50396 48372 50448
rect 50988 50396 51040 50448
rect 85856 50396 85908 50448
rect 90364 50396 90416 50448
rect 119436 50532 119488 50584
rect 119988 50532 120040 50584
rect 145840 50532 145892 50584
rect 146944 50532 146996 50584
rect 152924 50532 152976 50584
rect 168196 50532 168248 50584
rect 169668 50532 169720 50584
rect 188528 50532 188580 50584
rect 188988 50532 189040 50584
rect 204720 50532 204772 50584
rect 206928 50532 206980 50584
rect 219992 50532 220044 50584
rect 220728 50532 220780 50584
rect 232136 50532 232188 50584
rect 233148 50532 233200 50584
rect 242348 50532 242400 50584
rect 242808 50532 242860 50584
rect 250444 50532 250496 50584
rect 267004 50532 267056 50584
rect 270776 50532 270828 50584
rect 286968 50532 287020 50584
rect 289084 50532 289136 50584
rect 495256 50532 495308 50584
rect 504364 50532 504416 50584
rect 519636 50532 519688 50584
rect 554780 50532 554832 50584
rect 94044 50464 94096 50516
rect 118424 50464 118476 50516
rect 121368 50464 121420 50516
rect 146852 50464 146904 50516
rect 148968 50464 149020 50516
rect 170220 50464 170272 50516
rect 171048 50464 171100 50516
rect 189540 50464 189592 50516
rect 194508 50464 194560 50516
rect 209780 50464 209832 50516
rect 210976 50464 211028 50516
rect 224040 50464 224092 50516
rect 224868 50464 224920 50516
rect 235264 50464 235316 50516
rect 235816 50464 235868 50516
rect 245384 50464 245436 50516
rect 245568 50464 245620 50516
rect 253480 50464 253532 50516
rect 255228 50464 255280 50516
rect 261668 50464 261720 50516
rect 494244 50464 494296 50516
rect 515404 50464 515456 50516
rect 539600 50464 539652 50516
rect 568580 50464 568632 50516
rect 92388 50396 92440 50448
rect 121460 50396 121512 50448
rect 122748 50396 122800 50448
rect 147864 50396 147916 50448
rect 153016 50396 153068 50448
rect 174268 50396 174320 50448
rect 177856 50396 177908 50448
rect 194600 50396 194652 50448
rect 197268 50396 197320 50448
rect 211896 50396 211948 50448
rect 212448 50396 212500 50448
rect 225052 50396 225104 50448
rect 227536 50396 227588 50448
rect 238300 50396 238352 50448
rect 238668 50396 238720 50448
rect 247408 50396 247460 50448
rect 248328 50396 248380 50448
rect 255504 50396 255556 50448
rect 257988 50396 258040 50448
rect 263692 50396 263744 50448
rect 488172 50396 488224 50448
rect 497464 50396 497516 50448
rect 498384 50396 498436 50448
rect 525064 50396 525116 50448
rect 537944 50396 537996 50448
rect 575480 50396 575532 50448
rect 4068 50328 4120 50380
rect 46296 50328 46348 50380
rect 49608 50328 49660 50380
rect 84844 50328 84896 50380
rect 88248 50328 88300 50380
rect 124496 50328 124548 50380
rect 131580 50328 131632 50380
rect 132408 50328 132460 50380
rect 155960 50328 156012 50380
rect 158628 50328 158680 50380
rect 178316 50328 178368 50380
rect 179328 50328 179380 50380
rect 196624 50328 196676 50380
rect 202788 50328 202840 50380
rect 216956 50328 217008 50380
rect 217968 50328 218020 50380
rect 229100 50328 229152 50380
rect 230388 50328 230440 50380
rect 240324 50328 240376 50380
rect 244096 50328 244148 50380
rect 251456 50328 251508 50380
rect 252468 50328 252520 50380
rect 258632 50328 258684 50380
rect 277216 50328 277268 50380
rect 280896 50328 280948 50380
rect 343916 50328 343968 50380
rect 349252 50328 349304 50380
rect 440424 50328 440476 50380
rect 446404 50328 446456 50380
rect 474004 50328 474056 50380
rect 493324 50328 493376 50380
rect 503444 50328 503496 50380
rect 530584 50328 530636 50380
rect 534908 50328 534960 50380
rect 572812 50328 572864 50380
rect 33048 50260 33100 50312
rect 70676 50260 70728 50312
rect 75828 50260 75880 50312
rect 107200 50260 107252 50312
rect 111708 50260 111760 50312
rect 137652 50260 137704 50312
rect 143448 50260 143500 50312
rect 165160 50260 165212 50312
rect 169576 50260 169628 50312
rect 187516 50260 187568 50312
rect 191748 50260 191800 50312
rect 206744 50260 206796 50312
rect 209688 50260 209740 50312
rect 222016 50260 222068 50312
rect 527824 50260 527876 50312
rect 540244 50260 540296 50312
rect 28908 50192 28960 50244
rect 64144 50192 64196 50244
rect 26148 50124 26200 50176
rect 64512 50124 64564 50176
rect 74448 50192 74500 50244
rect 106188 50192 106240 50244
rect 106280 50192 106332 50244
rect 133604 50192 133656 50244
rect 134524 50192 134576 50244
rect 135628 50192 135680 50244
rect 142068 50192 142120 50244
rect 163780 50192 163832 50244
rect 164148 50192 164200 50244
rect 183376 50192 183428 50244
rect 184848 50192 184900 50244
rect 200672 50192 200724 50244
rect 201408 50192 201460 50244
rect 214932 50192 214984 50244
rect 531872 50192 531924 50244
rect 88892 50124 88944 50176
rect 113272 50124 113324 50176
rect 117228 50124 117280 50176
rect 142804 50124 142856 50176
rect 150348 50124 150400 50176
rect 171232 50124 171284 50176
rect 175188 50124 175240 50176
rect 192576 50124 192628 50176
rect 195888 50124 195940 50176
rect 210884 50124 210936 50176
rect 533896 50124 533948 50176
rect 545764 50124 545816 50176
rect 35808 50056 35860 50108
rect 72700 50056 72752 50108
rect 39948 49988 40000 50040
rect 76748 50056 76800 50108
rect 78588 50056 78640 50108
rect 85488 50056 85540 50108
rect 115388 50056 115440 50108
rect 118608 50056 118660 50108
rect 143816 50056 143868 50108
rect 147588 50056 147640 50108
rect 169208 50056 169260 50108
rect 176568 50056 176620 50108
rect 193588 50056 193640 50108
rect 83464 49988 83516 50040
rect 116400 49988 116452 50040
rect 45468 49920 45520 49972
rect 80796 49920 80848 49972
rect 82084 49920 82136 49972
rect 110236 49920 110288 49972
rect 119896 49920 119948 49972
rect 43444 49852 43496 49904
rect 69664 49852 69716 49904
rect 71136 49852 71188 49904
rect 73712 49852 73764 49904
rect 75184 49852 75236 49904
rect 104164 49852 104216 49904
rect 106924 49852 106976 49904
rect 125508 49988 125560 50040
rect 149888 49988 149940 50040
rect 154488 49988 154540 50040
rect 175280 49988 175332 50040
rect 177948 49988 178000 50040
rect 195612 49988 195664 50040
rect 263508 49988 263560 50040
rect 268752 49988 268804 50040
rect 144828 49920 144880 49972
rect 151728 49920 151780 49972
rect 172244 49920 172296 49972
rect 44824 49784 44876 49836
rect 60464 49784 60516 49836
rect 64236 49784 64288 49836
rect 46204 49716 46256 49768
rect 47308 49716 47360 49768
rect 50344 49716 50396 49768
rect 75736 49716 75788 49768
rect 76564 49716 76616 49768
rect 82820 49716 82872 49768
rect 86868 49784 86920 49836
rect 95884 49784 95936 49836
rect 122472 49784 122524 49836
rect 92020 49716 92072 49768
rect 93124 49716 93176 49768
rect 98092 49716 98144 49768
rect 98644 49716 98696 49768
rect 125140 49852 125192 49904
rect 124128 49784 124180 49836
rect 124864 49716 124916 49768
rect 140780 49852 140832 49904
rect 146208 49852 146260 49904
rect 153108 49852 153160 49904
rect 173256 49852 173308 49904
rect 173808 49920 173860 49972
rect 191564 49920 191616 49972
rect 193128 49920 193180 49972
rect 207756 49920 207808 49972
rect 270408 49920 270460 49972
rect 274824 49920 274876 49972
rect 177304 49852 177356 49904
rect 182088 49852 182140 49904
rect 198372 49852 198424 49904
rect 260656 49852 260708 49904
rect 266728 49852 266780 49904
rect 269028 49852 269080 49904
rect 273812 49852 273864 49904
rect 280068 49852 280120 49904
rect 283012 49852 283064 49904
rect 313464 49852 313516 49904
rect 314476 49852 314528 49904
rect 513564 49852 513616 49904
rect 519544 49852 519596 49904
rect 540980 49852 541032 49904
rect 548616 49852 548668 49904
rect 148876 49784 148928 49836
rect 155868 49784 155920 49836
rect 176292 49784 176344 49836
rect 249708 49784 249760 49836
rect 256516 49784 256568 49836
rect 259368 49784 259420 49836
rect 264704 49784 264756 49836
rect 271788 49784 271840 49836
rect 275836 49784 275888 49836
rect 281448 49784 281500 49836
rect 284024 49784 284076 49836
rect 288348 49784 288400 49836
rect 290096 49784 290148 49836
rect 317512 49784 317564 49836
rect 318708 49784 318760 49836
rect 319536 49784 319588 49836
rect 320824 49784 320876 49836
rect 336832 49784 336884 49836
rect 338856 49784 338908 49836
rect 434352 49784 434404 49836
rect 435364 49784 435416 49836
rect 451648 49784 451700 49836
rect 454684 49784 454736 49836
rect 137284 49716 137336 49768
rect 138756 49716 138808 49768
rect 157248 49716 157300 49768
rect 172428 49716 172480 49768
rect 251088 49716 251140 49768
rect 257528 49716 257580 49768
rect 260748 49716 260800 49768
rect 265716 49716 265768 49768
rect 268936 49716 268988 49768
rect 272800 49716 272852 49768
rect 273904 49716 273956 49768
rect 276848 49716 276900 49768
rect 278688 49716 278740 49768
rect 282000 49716 282052 49768
rect 282828 49716 282880 49768
rect 285036 49716 285088 49768
rect 289728 49716 289780 49768
rect 291108 49716 291160 49768
rect 312452 49716 312504 49768
rect 313464 49716 313516 49768
rect 316500 49716 316552 49768
rect 317604 49716 317656 49768
rect 320548 49716 320600 49768
rect 321468 49716 321520 49768
rect 321560 49716 321612 49768
rect 322756 49716 322808 49768
rect 324596 49716 324648 49768
rect 325516 49716 325568 49768
rect 328644 49716 328696 49768
rect 329748 49716 329800 49768
rect 331772 49716 331824 49768
rect 332508 49716 332560 49768
rect 333796 49716 333848 49768
rect 334624 49716 334676 49768
rect 335820 49716 335872 49768
rect 336648 49716 336700 49768
rect 337844 49716 337896 49768
rect 338764 49716 338816 49768
rect 339868 49716 339920 49768
rect 340788 49716 340840 49768
rect 340880 49716 340932 49768
rect 342168 49716 342220 49768
rect 347964 49716 348016 49768
rect 348976 49716 349028 49768
rect 351000 49716 351052 49768
rect 351828 49716 351880 49768
rect 352012 49716 352064 49768
rect 353116 49716 353168 49768
rect 355140 49716 355192 49768
rect 355968 49716 356020 49768
rect 356152 49716 356204 49768
rect 357348 49716 357400 49768
rect 359188 49716 359240 49768
rect 360108 49716 360160 49768
rect 360200 49716 360252 49768
rect 361488 49716 361540 49768
rect 363236 49716 363288 49768
rect 364156 49716 364208 49768
rect 367284 49716 367336 49768
rect 368296 49716 368348 49768
rect 370320 49716 370372 49768
rect 371148 49716 371200 49768
rect 371332 49716 371384 49768
rect 372528 49716 372580 49768
rect 374368 49716 374420 49768
rect 375288 49716 375340 49768
rect 375380 49716 375432 49768
rect 376576 49716 376628 49768
rect 378508 49716 378560 49768
rect 379428 49716 379480 49768
rect 379520 49716 379572 49768
rect 380716 49716 380768 49768
rect 382556 49716 382608 49768
rect 383476 49716 383528 49768
rect 386604 49716 386656 49768
rect 387708 49716 387760 49768
rect 389640 49716 389692 49768
rect 390468 49716 390520 49768
rect 390652 49716 390704 49768
rect 391756 49716 391808 49768
rect 393688 49716 393740 49768
rect 394608 49716 394660 49768
rect 394700 49716 394752 49768
rect 395896 49716 395948 49768
rect 397736 49716 397788 49768
rect 398656 49716 398708 49768
rect 400772 49716 400824 49768
rect 401508 49716 401560 49768
rect 401876 49716 401928 49768
rect 402888 49716 402940 49768
rect 405924 49716 405976 49768
rect 406936 49716 406988 49768
rect 408960 49716 409012 49768
rect 409788 49716 409840 49768
rect 409972 49716 410024 49768
rect 411076 49716 411128 49768
rect 413008 49716 413060 49768
rect 413928 49716 413980 49768
rect 414020 49716 414072 49768
rect 415308 49716 415360 49768
rect 417056 49716 417108 49768
rect 418068 49716 418120 49768
rect 420092 49716 420144 49768
rect 420828 49716 420880 49768
rect 421104 49716 421156 49768
rect 422208 49716 422260 49768
rect 424140 49716 424192 49768
rect 424968 49716 425020 49768
rect 425244 49716 425296 49768
rect 426256 49716 426308 49768
rect 428280 49716 428332 49768
rect 429108 49716 429160 49768
rect 429292 49716 429344 49768
rect 430488 49716 430540 49768
rect 432328 49716 432380 49768
rect 433248 49716 433300 49768
rect 433340 49716 433392 49768
rect 434628 49716 434680 49768
rect 436376 49716 436428 49768
rect 437388 49716 437440 49768
rect 439412 49716 439464 49768
rect 440148 49716 440200 49768
rect 443460 49716 443512 49768
rect 444288 49716 444340 49768
rect 444472 49716 444524 49768
rect 445668 49716 445720 49768
rect 447508 49716 447560 49768
rect 448428 49716 448480 49768
rect 448520 49716 448572 49768
rect 449808 49716 449860 49768
rect 452660 49716 452712 49768
rect 453856 49716 453908 49768
rect 455696 49716 455748 49768
rect 457444 49716 457496 49768
rect 459744 49716 459796 49768
rect 460756 49716 460808 49768
rect 462780 49716 462832 49768
rect 463608 49716 463660 49768
rect 463792 49716 463844 49768
rect 464988 49716 465040 49768
rect 466828 49716 466880 49768
rect 467748 49716 467800 49768
rect 467840 49716 467892 49768
rect 469036 49716 469088 49768
rect 470876 49716 470928 49768
rect 471796 49716 471848 49768
rect 475016 49716 475068 49768
rect 475936 49716 475988 49768
rect 478052 49716 478104 49768
rect 478788 49716 478840 49768
rect 479064 49716 479116 49768
rect 480168 49716 480220 49768
rect 482100 49716 482152 49768
rect 482928 49716 482980 49768
rect 483112 49716 483164 49768
rect 484216 49716 484268 49768
rect 486148 49716 486200 49768
rect 487068 49716 487120 49768
rect 487160 49716 487212 49768
rect 488448 49716 488500 49768
rect 490196 49716 490248 49768
rect 491116 49716 491168 49768
rect 497372 49716 497424 49768
rect 498108 49716 498160 49768
rect 501420 49716 501472 49768
rect 502248 49716 502300 49768
rect 502432 49716 502484 49768
rect 503628 49716 503680 49768
rect 505468 49716 505520 49768
rect 506388 49716 506440 49768
rect 517612 49716 517664 49768
rect 518716 49716 518768 49768
rect 520740 49716 520792 49768
rect 521568 49716 521620 49768
rect 521752 49716 521804 49768
rect 522948 49716 523000 49768
rect 524788 49716 524840 49768
rect 525708 49716 525760 49768
rect 532884 49716 532936 49768
rect 533988 49716 534040 49768
rect 535920 49716 535972 49768
rect 536748 49716 536800 49768
rect 536932 49716 536984 49768
rect 538128 49716 538180 49768
rect 539968 49716 540020 49768
rect 547144 49716 547196 49768
rect 66168 49580 66220 49632
rect 99104 49580 99156 49632
rect 70216 49512 70268 49564
rect 102140 49512 102192 49564
rect 41328 49444 41380 49496
rect 77208 49444 77260 49496
rect 84108 49444 84160 49496
rect 114284 49444 114336 49496
rect 34428 49376 34480 49428
rect 71688 49376 71740 49428
rect 73068 49376 73120 49428
rect 105176 49376 105228 49428
rect 7564 49308 7616 49360
rect 44272 49308 44324 49360
rect 52368 49308 52420 49360
rect 86500 49308 86552 49360
rect 102048 49308 102100 49360
rect 129556 49308 129608 49360
rect 298100 49308 298152 49360
rect 298836 49308 298888 49360
rect 37188 49240 37240 49292
rect 74724 49240 74776 49292
rect 79968 49240 80020 49292
rect 111248 49240 111300 49292
rect 129004 49240 129056 49292
rect 151912 49240 151964 49292
rect 4804 49172 4856 49224
rect 43260 49172 43312 49224
rect 48228 49172 48280 49224
rect 83832 49172 83884 49224
rect 86776 49172 86828 49224
rect 117412 49172 117464 49224
rect 131028 49172 131080 49224
rect 154948 49172 155000 49224
rect 17868 49104 17920 49156
rect 57428 49104 57480 49156
rect 62028 49104 62080 49156
rect 96068 49104 96120 49156
rect 97908 49104 97960 49156
rect 126520 49104 126572 49156
rect 129648 49104 129700 49156
rect 153936 49104 153988 49156
rect 8208 49036 8260 49088
rect 49332 49036 49384 49088
rect 59268 49036 59320 49088
rect 93032 49036 93084 49088
rect 104808 49036 104860 49088
rect 132592 49036 132644 49088
rect 133788 49036 133840 49088
rect 156972 49036 157024 49088
rect 3976 48968 4028 49020
rect 45284 48968 45336 49020
rect 55128 48968 55180 49020
rect 89904 48968 89956 49020
rect 91008 48968 91060 49020
rect 120448 48968 120500 49020
rect 126888 48968 126940 49020
rect 150900 48968 150952 49020
rect 555424 46860 555476 46912
rect 580172 46860 580224 46912
rect 293960 46112 294012 46164
rect 294788 46112 294840 46164
rect 3424 45500 3476 45552
rect 18604 45500 18656 45552
rect 3516 33056 3568 33108
rect 35164 33056 35216 33108
rect 574744 33056 574796 33108
rect 580172 33056 580224 33108
rect 108948 22720 109000 22772
rect 134524 22720 134576 22772
rect 30288 21360 30340 21412
rect 67732 21360 67784 21412
rect 3424 20612 3476 20664
rect 29644 20612 29696 20664
rect 566464 20612 566516 20664
rect 579988 20612 580040 20664
rect 151084 10276 151136 10328
rect 158812 10276 158864 10328
rect 3424 6808 3476 6860
rect 21364 6808 21416 6860
rect 551284 6808 551336 6860
rect 580172 6808 580224 6860
rect 21824 6128 21876 6180
rect 60740 6128 60792 6180
rect 520924 6128 520976 6180
rect 551468 6128 551520 6180
rect 556804 5516 556856 5568
rect 558552 5516 558604 5568
rect 560944 5516 560996 5568
rect 562048 5516 562100 5568
rect 504364 5380 504416 5432
rect 526628 5380 526680 5432
rect 500224 5312 500276 5364
rect 523040 5312 523092 5364
rect 482284 5244 482336 5296
rect 505376 5244 505428 5296
rect 461584 5176 461636 5228
rect 484032 5176 484084 5228
rect 487068 5176 487120 5228
rect 515956 5176 516008 5228
rect 446404 5108 446456 5160
rect 462780 5108 462832 5160
rect 480076 5108 480128 5160
rect 508872 5108 508924 5160
rect 462228 5040 462280 5092
rect 487620 5040 487672 5092
rect 489828 5040 489880 5092
rect 519452 5040 519504 5092
rect 519544 5040 519596 5092
rect 547880 5040 547932 5092
rect 431868 4972 431920 5024
rect 452108 4972 452160 5024
rect 464896 4972 464948 5024
rect 491024 4972 491076 5024
rect 502248 4972 502300 5024
rect 533712 4972 533764 5024
rect 536104 4972 536156 5024
rect 544384 4972 544436 5024
rect 429108 4904 429160 4956
rect 448612 4904 448664 4956
rect 469036 4904 469088 4956
rect 494704 4904 494756 4956
rect 505008 4904 505060 4956
rect 537208 4904 537260 4956
rect 93952 4836 94004 4888
rect 122840 4836 122892 4888
rect 437296 4836 437348 4888
rect 459192 4836 459244 4888
rect 471796 4836 471848 4888
rect 498200 4836 498252 4888
rect 507768 4836 507820 4888
rect 540796 4836 540848 4888
rect 76196 4768 76248 4820
rect 107660 4768 107712 4820
rect 435364 4768 435416 4820
rect 455696 4768 455748 4820
rect 457444 4768 457496 4820
rect 480536 4768 480588 4820
rect 484216 4768 484268 4820
rect 512460 4768 512512 4820
rect 518716 4768 518768 4820
rect 552664 4768 552716 4820
rect 62120 4632 62172 4684
rect 64880 4632 64932 4684
rect 525064 4632 525116 4684
rect 530124 4632 530176 4684
rect 51080 4496 51132 4548
rect 52460 4496 52512 4548
rect 493324 4428 493376 4480
rect 501788 4428 501840 4480
rect 38384 4088 38436 4140
rect 50344 4088 50396 4140
rect 342168 4088 342220 4140
rect 346952 4088 347004 4140
rect 348976 4088 349028 4140
rect 355232 4088 355284 4140
rect 365628 4088 365680 4140
rect 375288 4088 375340 4140
rect 378048 4088 378100 4140
rect 389456 4088 389508 4140
rect 397368 4088 397420 4140
rect 411904 4088 411956 4140
rect 415308 4088 415360 4140
rect 432052 4088 432104 4140
rect 433248 4088 433300 4140
rect 453304 4088 453356 4140
rect 460388 4088 460440 4140
rect 460756 4088 460808 4140
rect 485228 4088 485280 4140
rect 485688 4088 485740 4140
rect 514760 4088 514812 4140
rect 515404 4088 515456 4140
rect 525432 4088 525484 4140
rect 525708 4088 525760 4140
rect 560852 4088 560904 4140
rect 1676 4020 1728 4072
rect 7564 4020 7616 4072
rect 41880 4020 41932 4072
rect 53656 4020 53708 4072
rect 64144 4020 64196 4072
rect 314568 4020 314620 4072
rect 316224 4020 316276 4072
rect 332508 4020 332560 4072
rect 336280 4020 336332 4072
rect 340788 4020 340840 4072
rect 345756 4020 345808 4072
rect 351828 4020 351880 4072
rect 358728 4020 358780 4072
rect 367008 4020 367060 4072
rect 376484 4020 376536 4072
rect 382188 4020 382240 4072
rect 394240 4020 394292 4072
rect 395988 4020 396040 4072
rect 410800 4020 410852 4072
rect 411168 4020 411220 4072
rect 428464 4020 428516 4072
rect 430396 4020 430448 4072
rect 450912 4020 450964 4072
rect 456708 4020 456760 4072
rect 481732 4020 481784 4072
rect 484308 4020 484360 4072
rect 513564 4020 513616 4072
rect 518808 4020 518860 4072
rect 548616 4020 548668 4072
rect 549168 4020 549220 4072
rect 31300 3952 31352 4004
rect 43444 3952 43496 4004
rect 45376 3952 45428 4004
rect 71044 3952 71096 4004
rect 92756 3952 92808 4004
rect 95884 3952 95936 4004
rect 357348 3952 357400 4004
rect 364616 3952 364668 4004
rect 372528 3952 372580 4004
rect 382372 3952 382424 4004
rect 383476 3952 383528 4004
rect 395344 3952 395396 4004
rect 398656 3952 398708 4004
rect 413100 3952 413152 4004
rect 415216 3952 415268 4004
rect 433248 3952 433300 4004
rect 436008 3952 436060 4004
rect 456892 3952 456944 4004
rect 463608 3952 463660 4004
rect 488816 3952 488868 4004
rect 493968 3952 494020 4004
rect 524236 3952 524288 4004
rect 524328 3952 524380 4004
rect 559748 3952 559800 4004
rect 28816 3884 28868 3936
rect 55864 3884 55916 3936
rect 71504 3884 71556 3936
rect 75184 3884 75236 3936
rect 353208 3884 353260 3936
rect 361120 3884 361172 3936
rect 362868 3884 362920 3936
rect 371700 3884 371752 3936
rect 373908 3884 373960 3936
rect 384764 3884 384816 3936
rect 384948 3884 385000 3936
rect 397736 3884 397788 3936
rect 400128 3884 400180 3936
rect 415492 3884 415544 3936
rect 419448 3884 419500 3936
rect 437940 3884 437992 3936
rect 438768 3884 438820 3936
rect 453948 3884 454000 3936
rect 460848 3884 460900 3936
rect 486424 3884 486476 3936
rect 491116 3884 491168 3936
rect 520740 3884 520792 3936
rect 521568 3884 521620 3936
rect 553768 3884 553820 3936
rect 24216 3816 24268 3868
rect 54484 3816 54536 3868
rect 353116 3816 353168 3868
rect 359924 3816 359976 3868
rect 360108 3816 360160 3868
rect 368204 3816 368256 3868
rect 371148 3816 371200 3868
rect 381176 3816 381228 3868
rect 386328 3816 386380 3868
rect 398932 3816 398984 3868
rect 405648 3816 405700 3868
rect 421380 3816 421432 3868
rect 424968 3816 425020 3868
rect 443828 3816 443880 3868
rect 448428 3816 448480 3868
rect 471060 3816 471112 3868
rect 471888 3816 471940 3868
rect 499396 3816 499448 3868
rect 500868 3816 500920 3868
rect 532516 3816 532568 3868
rect 538128 3816 538180 3868
rect 575112 3816 575164 3868
rect 20536 3748 20588 3800
rect 44824 3748 44876 3800
rect 46664 3748 46716 3800
rect 76564 3748 76616 3800
rect 344928 3748 344980 3800
rect 351644 3748 351696 3800
rect 358636 3748 358688 3800
rect 367008 3748 367060 3800
rect 368296 3748 368348 3800
rect 377680 3748 377732 3800
rect 380808 3748 380860 3800
rect 393044 3748 393096 3800
rect 393228 3748 393280 3800
rect 407212 3748 407264 3800
rect 411076 3748 411128 3800
rect 427268 3748 427320 3800
rect 427728 3748 427780 3800
rect 447416 3748 447468 3800
rect 449808 3748 449860 3800
rect 472256 3748 472308 3800
rect 475936 3748 475988 3800
rect 502984 3748 503036 3800
rect 503628 3748 503680 3800
rect 534908 3748 534960 3800
rect 536748 3748 536800 3800
rect 573916 3748 573968 3800
rect 35992 3680 36044 3732
rect 71136 3680 71188 3732
rect 350448 3680 350500 3732
rect 357532 3680 357584 3732
rect 361488 3680 361540 3732
rect 369400 3680 369452 3732
rect 369768 3680 369820 3732
rect 379980 3680 380032 3732
rect 389088 3680 389140 3732
rect 402520 3680 402572 3732
rect 404268 3680 404320 3732
rect 420184 3680 420236 3732
rect 422208 3680 422260 3732
rect 440332 3680 440384 3732
rect 442908 3680 442960 3732
rect 465172 3680 465224 3732
rect 467748 3680 467800 3732
rect 493508 3680 493560 3732
rect 496728 3680 496780 3732
rect 527824 3680 527876 3732
rect 533988 3680 534040 3732
rect 570328 3680 570380 3732
rect 26516 3612 26568 3664
rect 572 3544 624 3596
rect 4804 3544 4856 3596
rect 12256 3544 12308 3596
rect 2872 3476 2924 3528
rect 3884 3476 3936 3528
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12348 3476 12400 3528
rect 15936 3544 15988 3596
rect 16488 3544 16540 3596
rect 17040 3544 17092 3596
rect 17868 3544 17920 3596
rect 18236 3544 18288 3596
rect 19248 3544 19300 3596
rect 19432 3544 19484 3596
rect 20628 3544 20680 3596
rect 25320 3544 25372 3596
rect 26148 3544 26200 3596
rect 27712 3544 27764 3596
rect 28908 3544 28960 3596
rect 32404 3544 32456 3596
rect 33048 3544 33100 3596
rect 33600 3544 33652 3596
rect 34428 3544 34480 3596
rect 43076 3612 43128 3664
rect 78864 3612 78916 3664
rect 96252 3612 96304 3664
rect 98644 3612 98696 3664
rect 62120 3544 62172 3596
rect 66720 3544 66772 3596
rect 67548 3544 67600 3596
rect 67916 3544 67968 3596
rect 68928 3544 68980 3596
rect 69112 3544 69164 3596
rect 70216 3544 70268 3596
rect 72608 3544 72660 3596
rect 73068 3544 73120 3596
rect 73804 3544 73856 3596
rect 74448 3544 74500 3596
rect 75000 3544 75052 3596
rect 75828 3544 75880 3596
rect 77392 3544 77444 3596
rect 78588 3544 78640 3596
rect 80888 3544 80940 3596
rect 81348 3544 81400 3596
rect 83280 3544 83332 3596
rect 84108 3544 84160 3596
rect 85672 3544 85724 3596
rect 86776 3544 86828 3596
rect 114008 3544 114060 3596
rect 124864 3544 124916 3596
rect 136456 3544 136508 3596
rect 151084 3612 151136 3664
rect 343548 3612 343600 3664
rect 349252 3612 349304 3664
rect 357256 3612 357308 3664
rect 365812 3612 365864 3664
rect 368388 3612 368440 3664
rect 378876 3612 378928 3664
rect 379428 3612 379480 3664
rect 390652 3612 390704 3664
rect 391756 3612 391808 3664
rect 404820 3612 404872 3664
rect 406936 3612 406988 3664
rect 422576 3612 422628 3664
rect 426256 3612 426308 3664
rect 445024 3612 445076 3664
rect 447048 3612 447100 3664
rect 469864 3612 469916 3664
rect 470508 3612 470560 3664
rect 497096 3612 497148 3664
rect 498108 3612 498160 3664
rect 529020 3612 529072 3664
rect 529848 3612 529900 3664
rect 566832 3612 566884 3664
rect 5264 3408 5316 3460
rect 46204 3408 46256 3460
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 44272 3340 44324 3392
rect 45468 3340 45520 3392
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 51356 3476 51408 3528
rect 52368 3476 52420 3528
rect 52552 3476 52604 3528
rect 53748 3476 53800 3528
rect 57152 3476 57204 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 60832 3476 60884 3528
rect 56048 3408 56100 3460
rect 56508 3408 56560 3460
rect 64328 3408 64380 3460
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 89168 3476 89220 3528
rect 90272 3476 90324 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 92388 3476 92440 3528
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 101036 3476 101088 3528
rect 102048 3476 102100 3528
rect 102232 3476 102284 3528
rect 103428 3476 103480 3528
rect 105728 3476 105780 3528
rect 106188 3476 106240 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 109316 3476 109368 3528
rect 110328 3476 110380 3528
rect 110512 3476 110564 3528
rect 111708 3476 111760 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 116400 3476 116452 3528
rect 117228 3476 117280 3528
rect 117596 3476 117648 3528
rect 118608 3476 118660 3528
rect 118792 3476 118844 3528
rect 119804 3476 119856 3528
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 125876 3476 125928 3528
rect 126888 3476 126940 3528
rect 126980 3476 127032 3528
rect 129004 3476 129056 3528
rect 130568 3476 130620 3528
rect 131028 3476 131080 3528
rect 146944 3544 146996 3596
rect 267740 3544 267792 3596
rect 268936 3544 268988 3596
rect 324228 3544 324280 3596
rect 326804 3544 326856 3596
rect 328368 3544 328420 3596
rect 331588 3544 331640 3596
rect 334624 3544 334676 3596
rect 338672 3544 338724 3596
rect 339408 3544 339460 3596
rect 344560 3544 344612 3596
rect 354588 3544 354640 3596
rect 362316 3544 362368 3596
rect 364156 3544 364208 3596
rect 372896 3544 372948 3596
rect 376576 3544 376628 3596
rect 387156 3544 387208 3596
rect 387616 3544 387668 3596
rect 401324 3544 401376 3596
rect 402796 3544 402848 3596
rect 418988 3544 419040 3596
rect 422116 3544 422168 3596
rect 441528 3544 441580 3596
rect 441620 3544 441672 3596
rect 463976 3544 464028 3596
rect 464988 3544 465040 3596
rect 489920 3544 489972 3596
rect 491208 3544 491260 3596
rect 521844 3544 521896 3596
rect 527088 3544 527140 3596
rect 563244 3544 563296 3596
rect 51080 3340 51132 3392
rect 78588 3340 78640 3392
rect 81992 3340 82044 3392
rect 82084 3340 82136 3392
rect 83464 3340 83516 3392
rect 88984 3408 89036 3460
rect 103336 3408 103388 3460
rect 106832 3408 106884 3460
rect 111616 3408 111668 3460
rect 93124 3340 93176 3392
rect 128176 3408 128228 3460
rect 142436 3476 142488 3528
rect 143448 3476 143500 3528
rect 143540 3476 143592 3528
rect 144644 3476 144696 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 149520 3476 149572 3528
rect 150348 3476 150400 3528
rect 150624 3476 150676 3528
rect 151728 3476 151780 3528
rect 151820 3476 151872 3528
rect 153108 3476 153160 3528
rect 155408 3476 155460 3528
rect 155868 3476 155920 3528
rect 156604 3476 156656 3528
rect 157248 3476 157300 3528
rect 157800 3476 157852 3528
rect 158628 3476 158680 3528
rect 158904 3476 158956 3528
rect 160008 3476 160060 3528
rect 160100 3476 160152 3528
rect 161388 3476 161440 3528
rect 163688 3476 163740 3528
rect 164148 3476 164200 3528
rect 166080 3476 166132 3528
rect 166908 3476 166960 3528
rect 167184 3476 167236 3528
rect 168288 3476 168340 3528
rect 168380 3476 168432 3528
rect 169484 3476 169536 3528
rect 171968 3476 172020 3528
rect 172428 3476 172480 3528
rect 173164 3476 173216 3528
rect 173808 3476 173860 3528
rect 174268 3476 174320 3528
rect 175188 3476 175240 3528
rect 175464 3476 175516 3528
rect 176568 3476 176620 3528
rect 176660 3476 176712 3528
rect 177764 3476 177816 3528
rect 180248 3476 180300 3528
rect 180708 3476 180760 3528
rect 181444 3476 181496 3528
rect 182088 3476 182140 3528
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 184940 3476 184992 3528
rect 186228 3476 186280 3528
rect 188528 3476 188580 3528
rect 188988 3476 189040 3528
rect 190828 3476 190880 3528
rect 191748 3476 191800 3528
rect 192024 3476 192076 3528
rect 193128 3476 193180 3528
rect 193220 3476 193272 3528
rect 194324 3476 194376 3528
rect 197912 3476 197964 3528
rect 198648 3476 198700 3528
rect 199108 3476 199160 3528
rect 200028 3476 200080 3528
rect 205088 3476 205140 3528
rect 205548 3476 205600 3528
rect 206192 3476 206244 3528
rect 206928 3476 206980 3528
rect 207388 3476 207440 3528
rect 208308 3476 208360 3528
rect 209780 3476 209832 3528
rect 211068 3476 211120 3528
rect 213368 3476 213420 3528
rect 213828 3476 213880 3528
rect 214472 3476 214524 3528
rect 215208 3476 215260 3528
rect 215668 3476 215720 3528
rect 216588 3476 216640 3528
rect 216864 3476 216916 3528
rect 217968 3476 218020 3528
rect 218060 3476 218112 3528
rect 219164 3476 219216 3528
rect 222752 3476 222804 3528
rect 223488 3476 223540 3528
rect 223948 3476 224000 3528
rect 224868 3476 224920 3528
rect 226340 3476 226392 3528
rect 227628 3476 227680 3528
rect 229836 3476 229888 3528
rect 230388 3476 230440 3528
rect 231032 3476 231084 3528
rect 231768 3476 231820 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 234620 3476 234672 3528
rect 235908 3476 235960 3528
rect 238116 3476 238168 3528
rect 238668 3476 238720 3528
rect 239312 3476 239364 3528
rect 240048 3476 240100 3528
rect 240508 3476 240560 3528
rect 241428 3476 241480 3528
rect 242900 3476 242952 3528
rect 244004 3476 244056 3528
rect 247592 3476 247644 3528
rect 248328 3476 248380 3528
rect 249984 3476 250036 3528
rect 251088 3476 251140 3528
rect 251180 3476 251232 3528
rect 252468 3476 252520 3528
rect 254676 3476 254728 3528
rect 255228 3476 255280 3528
rect 255872 3476 255924 3528
rect 256608 3476 256660 3528
rect 257068 3476 257120 3528
rect 257988 3476 258040 3528
rect 258264 3476 258316 3528
rect 259368 3476 259420 3528
rect 259460 3476 259512 3528
rect 260748 3476 260800 3528
rect 262956 3476 263008 3528
rect 263508 3476 263560 3528
rect 264152 3476 264204 3528
rect 264888 3476 264940 3528
rect 266544 3476 266596 3528
rect 267648 3476 267700 3528
rect 273628 3476 273680 3528
rect 274548 3476 274600 3528
rect 274824 3476 274876 3528
rect 275928 3476 275980 3528
rect 280712 3476 280764 3528
rect 281448 3476 281500 3528
rect 281908 3476 281960 3528
rect 282828 3476 282880 3528
rect 284300 3476 284352 3528
rect 285588 3476 285640 3528
rect 287796 3476 287848 3528
rect 288348 3476 288400 3528
rect 288992 3476 289044 3528
rect 289728 3476 289780 3528
rect 290188 3476 290240 3528
rect 291292 3476 291344 3528
rect 291384 3476 291436 3528
rect 292488 3476 292540 3528
rect 292580 3476 292632 3528
rect 294052 3476 294104 3528
rect 296076 3476 296128 3528
rect 296628 3476 296680 3528
rect 302424 3476 302476 3528
rect 303160 3476 303212 3528
rect 307760 3476 307812 3528
rect 309048 3476 309100 3528
rect 310428 3476 310480 3528
rect 311440 3476 311492 3528
rect 311808 3476 311860 3528
rect 312636 3476 312688 3528
rect 314476 3476 314528 3528
rect 315028 3476 315080 3528
rect 318708 3476 318760 3528
rect 319720 3476 319772 3528
rect 322756 3476 322808 3528
rect 324412 3476 324464 3528
rect 329748 3476 329800 3528
rect 332692 3476 332744 3528
rect 335268 3476 335320 3528
rect 336004 3476 336056 3528
rect 337476 3476 337528 3528
rect 338764 3476 338816 3528
rect 343364 3476 343416 3528
rect 347688 3476 347740 3528
rect 354036 3476 354088 3528
rect 355968 3476 356020 3528
rect 363512 3476 363564 3528
rect 364248 3476 364300 3528
rect 374092 3476 374144 3528
rect 376668 3476 376720 3528
rect 388260 3476 388312 3528
rect 391848 3476 391900 3528
rect 406016 3476 406068 3528
rect 407028 3476 407080 3528
rect 423772 3476 423824 3528
rect 426348 3476 426400 3528
rect 446220 3476 446272 3528
rect 449716 3476 449768 3528
rect 473452 3476 473504 3528
rect 476028 3476 476080 3528
rect 504180 3476 504232 3528
rect 506388 3476 506440 3528
rect 538404 3476 538456 3528
rect 539508 3476 539560 3528
rect 577412 3476 577464 3528
rect 134156 3408 134208 3460
rect 135168 3408 135220 3460
rect 138848 3408 138900 3460
rect 139308 3408 139360 3460
rect 141240 3408 141292 3460
rect 142068 3408 142120 3460
rect 161296 3408 161348 3460
rect 180064 3408 180116 3460
rect 189724 3408 189776 3460
rect 190368 3408 190420 3460
rect 265348 3408 265400 3460
rect 267004 3408 267056 3460
rect 272432 3408 272484 3460
rect 273904 3408 273956 3460
rect 321468 3408 321520 3460
rect 323308 3408 323360 3460
rect 325608 3408 325660 3460
rect 329196 3408 329248 3460
rect 331128 3408 331180 3460
rect 335084 3408 335136 3460
rect 339868 3408 339920 3460
rect 342076 3408 342128 3460
rect 348056 3408 348108 3460
rect 361396 3408 361448 3460
rect 370596 3408 370648 3460
rect 372436 3408 372488 3460
rect 383568 3408 383620 3460
rect 383660 3408 383712 3460
rect 396540 3408 396592 3460
rect 398748 3408 398800 3460
rect 414296 3408 414348 3460
rect 417976 3408 418028 3460
rect 436744 3408 436796 3460
rect 445576 3408 445628 3460
rect 468668 3408 468720 3460
rect 469128 3408 469180 3460
rect 495900 3408 495952 3460
rect 499488 3408 499540 3460
rect 530584 3408 530636 3460
rect 536104 3408 536156 3460
rect 582196 3408 582248 3460
rect 137284 3340 137336 3392
rect 329656 3340 329708 3392
rect 333888 3340 333940 3392
rect 375196 3340 375248 3392
rect 385960 3340 386012 3392
rect 387708 3340 387760 3392
rect 400128 3340 400180 3392
rect 401508 3340 401560 3392
rect 416688 3340 416740 3392
rect 423588 3340 423640 3392
rect 442632 3340 442684 3392
rect 455328 3340 455380 3392
rect 57244 3272 57296 3324
rect 64236 3272 64288 3324
rect 122288 3272 122340 3324
rect 122748 3272 122800 3324
rect 131764 3272 131816 3324
rect 132408 3272 132460 3324
rect 196808 3272 196860 3324
rect 197268 3272 197320 3324
rect 221556 3272 221608 3324
rect 222108 3272 222160 3324
rect 271236 3272 271288 3324
rect 271788 3272 271840 3324
rect 276020 3272 276072 3324
rect 277308 3272 277360 3324
rect 279516 3272 279568 3324
rect 280068 3272 280120 3324
rect 305000 3272 305052 3324
rect 305552 3272 305604 3324
rect 325516 3272 325568 3324
rect 328000 3272 328052 3324
rect 338856 3272 338908 3324
rect 342168 3272 342220 3324
rect 380716 3272 380768 3324
rect 391848 3272 391900 3324
rect 395896 3272 395948 3324
rect 409604 3272 409656 3324
rect 412548 3272 412600 3324
rect 429660 3272 429712 3324
rect 434628 3272 434680 3324
rect 454500 3272 454552 3324
rect 457996 3272 458048 3324
rect 478144 3340 478196 3392
rect 478788 3340 478840 3392
rect 506480 3340 506532 3392
rect 511908 3340 511960 3392
rect 545488 3340 545540 3392
rect 548524 3340 548576 3392
rect 583392 3340 583444 3392
rect 132960 3204 133012 3256
rect 133788 3204 133840 3256
rect 183744 3204 183796 3256
rect 184848 3204 184900 3256
rect 200304 3204 200356 3256
rect 201408 3204 201460 3256
rect 225144 3204 225196 3256
rect 226248 3204 226300 3256
rect 309140 3204 309192 3256
rect 310244 3204 310296 3256
rect 322848 3204 322900 3256
rect 325608 3204 325660 3256
rect 336648 3204 336700 3256
rect 340972 3204 341024 3256
rect 402888 3204 402940 3256
rect 417884 3204 417936 3256
rect 418068 3204 418120 3256
rect 435548 3204 435600 3256
rect 437388 3204 437440 3256
rect 458088 3204 458140 3256
rect 479340 3272 479392 3324
rect 481548 3272 481600 3324
rect 510068 3272 510120 3324
rect 514668 3272 514720 3324
rect 549076 3272 549128 3324
rect 549168 3272 549220 3324
rect 581000 3272 581052 3324
rect 482836 3204 482888 3256
rect 488448 3204 488500 3256
rect 517152 3204 517204 3256
rect 522948 3204 523000 3256
rect 557356 3204 557408 3256
rect 241704 3136 241756 3188
rect 242808 3136 242860 3188
rect 283104 3136 283156 3188
rect 285772 3136 285824 3188
rect 326988 3136 327040 3188
rect 330392 3136 330444 3188
rect 390468 3136 390520 3188
rect 403624 3136 403676 3188
rect 408316 3136 408368 3188
rect 246396 3068 246448 3120
rect 246948 3068 247000 3120
rect 297272 3068 297324 3120
rect 298192 3068 298244 3120
rect 394608 3068 394660 3120
rect 408408 3068 408460 3120
rect 420828 3136 420880 3188
rect 439136 3136 439188 3188
rect 453856 3136 453908 3188
rect 476948 3136 477000 3188
rect 482928 3136 482980 3188
rect 511264 3136 511316 3188
rect 516048 3136 516100 3188
rect 550272 3136 550324 3188
rect 556160 3136 556212 3188
rect 424968 3068 425020 3120
rect 430488 3068 430540 3120
rect 449808 3068 449860 3120
rect 451188 3068 451240 3120
rect 474556 3068 474608 3120
rect 480168 3068 480220 3120
rect 507676 3068 507728 3120
rect 513288 3068 513340 3120
rect 546684 3068 546736 3120
rect 547144 3068 547196 3120
rect 578608 3068 578660 3120
rect 135260 3000 135312 3052
rect 136548 3000 136600 3052
rect 140044 3000 140096 3052
rect 140688 3000 140740 3052
rect 164884 3000 164936 3052
rect 165528 3000 165580 3052
rect 201500 3000 201552 3052
rect 202604 3000 202656 3052
rect 208584 3000 208636 3052
rect 209688 3000 209740 3052
rect 248788 3000 248840 3052
rect 249708 3000 249760 3052
rect 318616 3000 318668 3052
rect 320916 3000 320968 3052
rect 346308 3000 346360 3052
rect 352840 3000 352892 3052
rect 416596 3000 416648 3052
rect 434444 3000 434496 3052
rect 445668 3000 445720 3052
rect 467472 3000 467524 3052
rect 473268 3000 473320 3052
rect 500592 3000 500644 3052
rect 509148 3000 509200 3052
rect 541992 3000 542044 3052
rect 542268 3000 542320 3052
rect 571524 3000 571576 3052
rect 320824 2932 320876 2984
rect 322112 2932 322164 2984
rect 349068 2932 349120 2984
rect 356336 2932 356388 2984
rect 413928 2932 413980 2984
rect 430856 2932 430908 2984
rect 440148 2932 440200 2984
rect 461584 2932 461636 2984
rect 466368 2932 466420 2984
rect 492312 2932 492364 2984
rect 497464 2932 497516 2984
rect 518348 2932 518400 2984
rect 531320 2932 531372 2984
rect 540244 2932 540296 2984
rect 564440 2932 564492 2984
rect 65524 2864 65576 2916
rect 66168 2864 66220 2916
rect 409788 2864 409840 2916
rect 426164 2864 426216 2916
rect 444288 2864 444340 2916
rect 466276 2864 466328 2916
rect 545764 2864 545816 2916
rect 294880 2796 294932 2848
rect 295432 2796 295484 2848
rect 454684 2796 454736 2848
rect 475752 2796 475804 2848
rect 544476 2796 544528 2848
rect 568028 2864 568080 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700670 73016 703520
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 105464 699718 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 170324 699718 170352 703520
rect 202800 700126 202828 703520
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 218992 700058 219020 703520
rect 218980 700052 219032 700058
rect 218980 699994 219032 700000
rect 235184 699718 235212 703520
rect 260748 700868 260800 700874
rect 260748 700810 260800 700816
rect 246948 700596 247000 700602
rect 246948 700538 247000 700544
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 173164 699712 173216 699718
rect 173164 699654 173216 699660
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 240784 699712 240836 699718
rect 240784 699654 240836 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 106200 659054 106228 699654
rect 173176 659190 173204 699654
rect 234528 696992 234580 696998
rect 234528 696934 234580 696940
rect 229836 670812 229888 670818
rect 229836 670754 229888 670760
rect 173164 659184 173216 659190
rect 173164 659126 173216 659132
rect 106188 659048 106240 659054
rect 106188 658990 106240 658996
rect 29644 658368 29696 658374
rect 29644 658310 29696 658316
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 658102 3464 658135
rect 3424 658096 3476 658102
rect 3424 658038 3476 658044
rect 25596 657756 25648 657762
rect 25596 657698 25648 657704
rect 4802 657520 4858 657529
rect 4802 657455 4858 657464
rect 3422 654256 3478 654265
rect 3422 654191 3478 654200
rect 3332 633412 3384 633418
rect 3332 633354 3384 633360
rect 3344 632097 3372 633354
rect 3330 632088 3386 632097
rect 3330 632023 3386 632032
rect 3148 619336 3200 619342
rect 3148 619278 3200 619284
rect 3160 619177 3188 619278
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3056 607164 3108 607170
rect 3056 607106 3108 607112
rect 3068 606121 3096 607106
rect 3054 606112 3110 606121
rect 3054 606047 3110 606056
rect 3332 580984 3384 580990
rect 3332 580926 3384 580932
rect 3344 580009 3372 580926
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3332 567180 3384 567186
rect 3332 567122 3384 567128
rect 3344 566953 3372 567122
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3332 554736 3384 554742
rect 3332 554678 3384 554684
rect 3344 553897 3372 554678
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3332 528556 3384 528562
rect 3332 528498 3384 528504
rect 3344 527921 3372 528498
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3148 516112 3200 516118
rect 3148 516054 3200 516060
rect 3160 514865 3188 516054
rect 3146 514856 3202 514865
rect 3146 514791 3202 514800
rect 2964 502308 3016 502314
rect 2964 502250 3016 502256
rect 2976 501809 3004 502250
rect 2962 501800 3018 501809
rect 2962 501735 3018 501744
rect 3240 476060 3292 476066
rect 3240 476002 3292 476008
rect 3252 475697 3280 476002
rect 3238 475688 3294 475697
rect 3238 475623 3294 475632
rect 3056 463684 3108 463690
rect 3056 463626 3108 463632
rect 3068 462641 3096 463626
rect 3054 462632 3110 462641
rect 3054 462567 3110 462576
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3332 293956 3384 293962
rect 3332 293898 3384 293904
rect 3344 293185 3372 293898
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3332 215008 3384 215014
rect 3330 214976 3332 214985
rect 3384 214976 3386 214985
rect 3330 214911 3386 214920
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 97617 3464 654191
rect 3516 654152 3568 654158
rect 3516 654094 3568 654100
rect 3528 201929 3556 654094
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 4816 58682 4844 657455
rect 11704 657348 11756 657354
rect 11704 657290 11756 657296
rect 7564 655716 7616 655722
rect 7564 655658 7616 655664
rect 7576 215014 7604 655658
rect 7656 655172 7708 655178
rect 7656 655114 7708 655120
rect 7668 619342 7696 655114
rect 10324 655036 10376 655042
rect 10324 654978 10376 654984
rect 7656 619336 7708 619342
rect 7656 619278 7708 619284
rect 10336 567186 10364 654978
rect 10324 567180 10376 567186
rect 10324 567122 10376 567128
rect 11716 306338 11744 657290
rect 15844 657076 15896 657082
rect 15844 657018 15896 657024
rect 11888 656668 11940 656674
rect 11888 656610 11940 656616
rect 11796 654764 11848 654770
rect 11796 654706 11848 654712
rect 11808 398818 11836 654706
rect 11900 633418 11928 656610
rect 14556 656532 14608 656538
rect 14556 656474 14608 656480
rect 14464 654492 14516 654498
rect 14464 654434 14516 654440
rect 11888 633412 11940 633418
rect 11888 633354 11940 633360
rect 11796 398812 11848 398818
rect 11796 398754 11848 398760
rect 11704 306332 11756 306338
rect 11704 306274 11756 306280
rect 14476 293962 14504 654434
rect 14568 580990 14596 656474
rect 14556 580984 14608 580990
rect 14556 580926 14608 580932
rect 14464 293956 14516 293962
rect 14464 293898 14516 293904
rect 7564 215008 7616 215014
rect 7564 214950 7616 214956
rect 15856 189038 15884 657018
rect 15936 656464 15988 656470
rect 15936 656406 15988 656412
rect 15948 528562 15976 656406
rect 17316 656396 17368 656402
rect 17316 656338 17368 656344
rect 17222 654392 17278 654401
rect 17222 654327 17278 654336
rect 15936 528556 15988 528562
rect 15936 528498 15988 528504
rect 15844 189032 15896 189038
rect 15844 188974 15896 188980
rect 17236 85542 17264 654327
rect 17328 476066 17356 656338
rect 18696 656260 18748 656266
rect 18696 656202 18748 656208
rect 18602 653712 18658 653721
rect 18602 653647 18658 653656
rect 17316 476060 17368 476066
rect 17316 476002 17368 476008
rect 17224 85536 17276 85542
rect 17224 85478 17276 85484
rect 2780 58676 2832 58682
rect 2780 58618 2832 58624
rect 4804 58676 4856 58682
rect 4804 58618 4856 58624
rect 2792 58585 2820 58618
rect 2778 58576 2834 58585
rect 2778 58511 2834 58520
rect 16488 50924 16540 50930
rect 16488 50866 16540 50872
rect 12348 50856 12400 50862
rect 12348 50798 12400 50804
rect 10968 50720 11020 50726
rect 10968 50662 11020 50668
rect 9588 50516 9640 50522
rect 9588 50458 9640 50464
rect 6828 50448 6880 50454
rect 6828 50390 6880 50396
rect 4068 50380 4120 50386
rect 4068 50322 4120 50328
rect 3976 49020 4028 49026
rect 3976 48962 4028 48968
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3988 6914 4016 48962
rect 3896 6886 4016 6914
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 572 3596 624 3602
rect 572 3538 624 3544
rect 584 480 612 3538
rect 1688 480 1716 4014
rect 3896 3534 3924 6886
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 2884 480 2912 3470
rect 4080 480 4108 50322
rect 4804 49224 4856 49230
rect 4804 49166 4856 49172
rect 4816 3602 4844 49166
rect 6840 6914 6868 50390
rect 7564 49360 7616 49366
rect 7564 49302 7616 49308
rect 6472 6886 6868 6914
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6472 480 6500 6886
rect 7576 4078 7604 49302
rect 8208 49088 8260 49094
rect 8208 49030 8260 49036
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 8220 3534 8248 49030
rect 9600 3534 9628 50458
rect 10980 3534 11008 50662
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 7668 480 7696 3470
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 12268 1850 12296 3538
rect 12360 3534 12388 50798
rect 15108 50652 15160 50658
rect 15108 50594 15160 50600
rect 13728 50584 13780 50590
rect 13728 50526 13780 50532
rect 13740 6914 13768 50526
rect 15120 6914 15148 50594
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12268 1822 12388 1850
rect 12360 480 12388 1822
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3602 16528 50866
rect 17868 49156 17920 49162
rect 17868 49098 17920 49104
rect 17880 3602 17908 49098
rect 18616 45558 18644 653647
rect 18708 423638 18736 656202
rect 21456 656124 21508 656130
rect 21456 656066 21508 656072
rect 21362 653576 21418 653585
rect 21362 653511 21418 653520
rect 18696 423632 18748 423638
rect 18696 423574 18748 423580
rect 19248 50992 19300 50998
rect 19248 50934 19300 50940
rect 18604 45552 18656 45558
rect 18604 45494 18656 45500
rect 19260 3602 19288 50934
rect 20628 50788 20680 50794
rect 20628 50730 20680 50736
rect 20536 3800 20588 3806
rect 20536 3742 20588 3748
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 15948 480 15976 3538
rect 17052 480 17080 3538
rect 18248 480 18276 3538
rect 19444 480 19472 3538
rect 20548 1986 20576 3742
rect 20640 3602 20668 50730
rect 21376 6866 21404 653511
rect 21468 372570 21496 656066
rect 22744 656056 22796 656062
rect 22744 655998 22796 656004
rect 21456 372564 21508 372570
rect 21456 372506 21508 372512
rect 22756 320142 22784 655998
rect 25504 655988 25556 655994
rect 25504 655930 25556 655936
rect 22836 654968 22888 654974
rect 22836 654910 22888 654916
rect 22848 463690 22876 654910
rect 22836 463684 22888 463690
rect 22836 463626 22888 463632
rect 22744 320136 22796 320142
rect 22744 320078 22796 320084
rect 25516 267714 25544 655930
rect 25608 411262 25636 657698
rect 26884 654696 26936 654702
rect 26884 654638 26936 654644
rect 25596 411256 25648 411262
rect 25596 411198 25648 411204
rect 26896 358766 26924 654638
rect 26884 358760 26936 358766
rect 26884 358702 26936 358708
rect 25504 267708 25556 267714
rect 25504 267650 25556 267656
rect 23388 51060 23440 51066
rect 23388 51002 23440 51008
rect 23400 6914 23428 51002
rect 28908 50244 28960 50250
rect 28908 50186 28960 50192
rect 26148 50176 26200 50182
rect 26148 50118 26200 50124
rect 23032 6886 23428 6914
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20548 1958 20668 1986
rect 20640 480 20668 1958
rect 21836 480 21864 6122
rect 23032 480 23060 6886
rect 24216 3868 24268 3874
rect 24216 3810 24268 3816
rect 24228 480 24256 3810
rect 26160 3602 26188 50118
rect 28816 3936 28868 3942
rect 28816 3878 28868 3884
rect 26516 3664 26568 3670
rect 26516 3606 26568 3612
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 25332 480 25360 3538
rect 26528 480 26556 3606
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27724 480 27752 3538
rect 28828 1986 28856 3878
rect 28920 3602 28948 50186
rect 29656 20670 29684 658310
rect 53656 658300 53708 658306
rect 53656 658242 53708 658248
rect 42248 658028 42300 658034
rect 42248 657970 42300 657976
rect 39304 657484 39356 657490
rect 39304 657426 39356 657432
rect 36544 657416 36596 657422
rect 36544 657358 36596 657364
rect 33782 656024 33838 656033
rect 33782 655959 33838 655968
rect 29736 655852 29788 655858
rect 29736 655794 29788 655800
rect 29748 164218 29776 655794
rect 32404 655648 32456 655654
rect 32404 655590 32456 655596
rect 29736 164212 29788 164218
rect 29736 164154 29788 164160
rect 32416 111790 32444 655590
rect 32404 111784 32456 111790
rect 32404 111726 32456 111732
rect 33796 71738 33824 655959
rect 35162 655888 35218 655897
rect 35162 655823 35218 655832
rect 33784 71732 33836 71738
rect 33784 71674 33836 71680
rect 33048 50312 33100 50318
rect 33048 50254 33100 50260
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 29644 20664 29696 20670
rect 29644 20606 29696 20612
rect 30300 6914 30328 21354
rect 30116 6886 30328 6914
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28828 1958 28948 1986
rect 28920 480 28948 1958
rect 30116 480 30144 6886
rect 31300 4004 31352 4010
rect 31300 3946 31352 3952
rect 31312 480 31340 3946
rect 33060 3602 33088 50254
rect 34428 49428 34480 49434
rect 34428 49370 34480 49376
rect 34440 3602 34468 49370
rect 35176 33114 35204 655823
rect 36556 255270 36584 657358
rect 36636 654900 36688 654906
rect 36636 654842 36688 654848
rect 36648 346390 36676 654842
rect 36726 653304 36782 653313
rect 36726 653239 36782 653248
rect 36740 607170 36768 653239
rect 36728 607164 36780 607170
rect 36728 607106 36780 607112
rect 36636 346384 36688 346390
rect 36636 346326 36688 346332
rect 36544 255264 36596 255270
rect 36544 255206 36596 255212
rect 39316 241466 39344 657426
rect 42064 657212 42116 657218
rect 42064 657154 42116 657160
rect 40776 655240 40828 655246
rect 40776 655182 40828 655188
rect 40682 654664 40738 654673
rect 40682 654599 40738 654608
rect 39394 653984 39450 653993
rect 39394 653919 39450 653928
rect 39408 554742 39436 653919
rect 39396 554736 39448 554742
rect 39396 554678 39448 554684
rect 39304 241460 39356 241466
rect 39304 241402 39356 241408
rect 40696 137970 40724 654599
rect 40788 502314 40816 655182
rect 40776 502308 40828 502314
rect 40776 502250 40828 502256
rect 42076 150414 42104 657154
rect 42156 655104 42208 655110
rect 42156 655046 42208 655052
rect 42168 449886 42196 655046
rect 42260 516118 42288 657970
rect 45190 655616 45246 655625
rect 44942 655574 45190 655602
rect 53668 655588 53696 658242
rect 211804 658232 211856 658238
rect 211804 658174 211856 658180
rect 194232 658164 194284 658170
rect 194232 658106 194284 658112
rect 132776 657960 132828 657966
rect 132776 657902 132828 657908
rect 184848 657960 184900 657966
rect 184848 657902 184900 657908
rect 185492 657960 185544 657966
rect 185492 657902 185544 657908
rect 80058 657384 80114 657393
rect 80058 657319 80114 657328
rect 62486 657248 62542 657257
rect 62486 657183 62542 657192
rect 58438 655752 58494 655761
rect 58438 655687 58494 655696
rect 58452 655602 58480 655687
rect 58098 655574 58480 655602
rect 62500 655588 62528 657183
rect 66810 657112 66866 657121
rect 66810 657047 66866 657056
rect 66824 655588 66852 657047
rect 75644 657008 75696 657014
rect 75644 656950 75696 656956
rect 71254 655586 71544 655602
rect 75656 655588 75684 656950
rect 80072 655588 80100 657319
rect 110788 657280 110840 657286
rect 110788 657222 110840 657228
rect 88800 657144 88852 657150
rect 88800 657086 88852 657092
rect 84384 656940 84436 656946
rect 84384 656882 84436 656888
rect 84396 655588 84424 656882
rect 88812 655588 88840 657086
rect 97632 655784 97684 655790
rect 97632 655726 97684 655732
rect 97644 655588 97672 655726
rect 110800 655588 110828 657222
rect 123944 655920 123996 655926
rect 123944 655862 123996 655868
rect 123956 655588 123984 655862
rect 132788 655588 132816 657902
rect 167920 657892 167972 657898
rect 167920 657834 167972 657840
rect 163504 657688 163556 657694
rect 163504 657630 163556 657636
rect 154672 657620 154724 657626
rect 154672 657562 154724 657568
rect 137100 657552 137152 657558
rect 137100 657494 137152 657500
rect 137112 655588 137140 657494
rect 154684 655588 154712 657562
rect 159088 656328 159140 656334
rect 159088 656270 159140 656276
rect 159100 655588 159128 656270
rect 163516 655588 163544 657630
rect 167932 655588 167960 657834
rect 181076 657824 181128 657830
rect 181076 657766 181128 657772
rect 176660 656600 176712 656606
rect 176660 656542 176712 656548
rect 172244 656192 172296 656198
rect 172244 656134 172296 656140
rect 172256 655588 172284 656134
rect 176672 655588 176700 656542
rect 181088 655588 181116 657766
rect 71254 655580 71556 655586
rect 71254 655574 71504 655580
rect 45190 655551 45246 655560
rect 71504 655522 71556 655528
rect 184860 655450 184888 657902
rect 185504 655588 185532 657902
rect 189816 656736 189868 656742
rect 189816 656678 189868 656684
rect 189828 655588 189856 656678
rect 194244 655588 194272 658106
rect 203064 656804 203116 656810
rect 203064 656746 203116 656752
rect 203076 655588 203104 656746
rect 211816 655588 211844 658174
rect 216220 656872 216272 656878
rect 216220 656814 216272 656820
rect 216232 655588 216260 656814
rect 229848 655602 229876 670754
rect 234540 663794 234568 696934
rect 238668 683256 238720 683262
rect 238668 683198 238720 683204
rect 234264 663766 234568 663794
rect 234264 655602 234292 663766
rect 238680 655602 238708 683198
rect 240796 659326 240824 699654
rect 240784 659320 240836 659326
rect 240784 659262 240836 659268
rect 242532 658980 242584 658986
rect 242532 658922 242584 658928
rect 229402 655574 229876 655602
rect 233818 655574 234292 655602
rect 238234 655574 238708 655602
rect 242544 655588 242572 658922
rect 246960 655588 246988 700538
rect 252468 700528 252520 700534
rect 252468 700470 252520 700476
rect 252480 663794 252508 700470
rect 260760 663794 260788 700810
rect 264888 700800 264940 700806
rect 264888 700742 264940 700748
rect 251744 663766 252508 663794
rect 260576 663766 260788 663794
rect 251744 655602 251772 663766
rect 255780 659252 255832 659258
rect 255780 659194 255832 659200
rect 251390 655574 251772 655602
rect 255792 655588 255820 659194
rect 260576 655602 260604 663766
rect 264900 655602 264928 700742
rect 267660 699854 267688 703520
rect 278688 700256 278740 700262
rect 278688 700198 278740 700204
rect 274548 700188 274600 700194
rect 274548 700130 274600 700136
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 274560 663794 274588 700130
rect 278700 663794 278728 700198
rect 283852 699786 283880 703520
rect 291108 699984 291160 699990
rect 291108 699926 291160 699932
rect 286968 699916 287020 699922
rect 286968 699858 287020 699864
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 286980 663794 287008 699858
rect 273824 663766 274588 663794
rect 278056 663766 278728 663794
rect 286888 663766 287008 663794
rect 268936 659116 268988 659122
rect 268936 659058 268988 659064
rect 260130 655574 260604 655602
rect 264546 655574 264928 655602
rect 268948 655588 268976 659058
rect 273824 655602 273852 663766
rect 278056 655602 278084 663766
rect 282092 660340 282144 660346
rect 282092 660282 282144 660288
rect 273378 655574 273852 655602
rect 277702 655574 278084 655602
rect 282104 655588 282132 660282
rect 286888 655602 286916 663766
rect 291120 655602 291148 699926
rect 299572 699848 299624 699854
rect 299572 699790 299624 699796
rect 296628 698964 296680 698970
rect 296628 698906 296680 698912
rect 296640 663794 296668 698906
rect 295720 663766 296668 663794
rect 295720 655602 295748 663766
rect 286534 655574 286916 655602
rect 290950 655574 291148 655602
rect 295366 655574 295748 655602
rect 299584 655602 299612 699790
rect 300136 698970 300164 703520
rect 329840 701004 329892 701010
rect 329840 700946 329892 700952
rect 325700 700936 325752 700942
rect 325700 700878 325752 700884
rect 311900 700120 311952 700126
rect 311900 700062 311952 700068
rect 303620 699780 303672 699786
rect 303620 699722 303672 699728
rect 300124 698964 300176 698970
rect 300124 698906 300176 698912
rect 303632 673454 303660 699722
rect 311912 673454 311940 700062
rect 316040 700052 316092 700058
rect 316040 699994 316092 700000
rect 316052 673454 316080 699994
rect 303632 673426 303752 673454
rect 311912 673426 312584 673454
rect 316052 673426 316816 673454
rect 303724 655602 303752 673426
rect 308496 659320 308548 659326
rect 308496 659262 308548 659268
rect 299584 655574 299690 655602
rect 303724 655574 304106 655602
rect 308508 655588 308536 659262
rect 312556 655602 312584 673426
rect 316788 655602 316816 673426
rect 321652 659184 321704 659190
rect 321652 659126 321704 659132
rect 312556 655574 312938 655602
rect 316788 655574 317262 655602
rect 321664 655588 321692 659126
rect 325712 655602 325740 700878
rect 329852 673454 329880 700946
rect 332520 699922 332548 703520
rect 336004 700936 336056 700942
rect 336004 700878 336056 700884
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 329852 673426 330064 673454
rect 330036 655602 330064 673426
rect 336016 660346 336044 700878
rect 343640 700732 343692 700738
rect 343640 700674 343692 700680
rect 338120 700664 338172 700670
rect 338120 700606 338172 700612
rect 340144 700664 340196 700670
rect 340144 700606 340196 700612
rect 338132 673454 338160 700606
rect 338132 673426 338896 673454
rect 336004 660340 336056 660346
rect 336004 660282 336056 660288
rect 334808 659048 334860 659054
rect 334808 658990 334860 658996
rect 325712 655574 326094 655602
rect 330036 655574 330510 655602
rect 334820 655588 334848 658990
rect 338868 655602 338896 673426
rect 340156 659258 340184 700606
rect 340144 659252 340196 659258
rect 340144 659194 340196 659200
rect 338868 655574 339250 655602
rect 343652 655588 343680 700674
rect 347780 700460 347832 700466
rect 347780 700402 347832 700408
rect 347792 655602 347820 700402
rect 348804 699990 348832 703520
rect 364996 700942 365024 703520
rect 364984 700936 365036 700942
rect 364984 700878 365036 700884
rect 356060 700392 356112 700398
rect 356060 700334 356112 700340
rect 351920 700324 351972 700330
rect 351920 700266 351972 700272
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 351932 655602 351960 700266
rect 356072 673454 356100 700334
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 360200 683188 360252 683194
rect 360200 683130 360252 683136
rect 360212 673454 360240 683130
rect 356072 673426 356376 673454
rect 360212 673426 360792 673454
rect 356348 655602 356376 673426
rect 360764 655602 360792 673426
rect 369860 670744 369912 670750
rect 369860 670686 369912 670692
rect 365628 658096 365680 658102
rect 365628 658038 365680 658044
rect 347792 655574 348082 655602
rect 351932 655574 352406 655602
rect 356348 655574 356822 655602
rect 360764 655574 361238 655602
rect 365640 655588 365668 658038
rect 369872 655602 369900 670686
rect 429212 659122 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 494808 700670 494836 703520
rect 494796 700664 494848 700670
rect 494796 700606 494848 700612
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 559668 700330 559696 703520
rect 543004 700324 543056 700330
rect 543004 700266 543056 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 429200 659116 429252 659122
rect 429200 659058 429252 659064
rect 543016 658986 543044 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 543004 658980 543056 658986
rect 543004 658922 543056 658928
rect 541348 658368 541400 658374
rect 541348 658310 541400 658316
rect 409512 658028 409564 658034
rect 409512 657970 409564 657976
rect 374368 656668 374420 656674
rect 374368 656610 374420 656616
rect 369872 655574 369978 655602
rect 374380 655588 374408 656610
rect 387524 656532 387576 656538
rect 387524 656474 387576 656480
rect 387536 655588 387564 656474
rect 400772 656464 400824 656470
rect 400772 656406 400824 656412
rect 400784 655588 400812 656406
rect 409524 655588 409552 657970
rect 435916 657756 435968 657762
rect 435916 657698 435968 657704
rect 413928 656396 413980 656402
rect 413928 656338 413980 656344
rect 413940 655588 413968 656338
rect 427084 656260 427136 656266
rect 427084 656202 427136 656208
rect 427096 655588 427124 656202
rect 435928 655588 435956 657698
rect 528098 657520 528154 657529
rect 471060 657484 471112 657490
rect 528098 657455 528154 657464
rect 471060 657426 471112 657432
rect 462228 657348 462280 657354
rect 462228 657290 462280 657296
rect 440240 656124 440292 656130
rect 440240 656066 440292 656072
rect 440252 655588 440280 656066
rect 453488 656056 453540 656062
rect 453488 655998 453540 656004
rect 453500 655588 453528 655998
rect 462240 655588 462268 657290
rect 466644 655988 466696 655994
rect 466644 655930 466696 655936
rect 466656 655588 466684 655930
rect 471072 655588 471100 657426
rect 475384 657416 475436 657422
rect 475384 657358 475436 657364
rect 475396 655588 475424 657358
rect 501788 657212 501840 657218
rect 501788 657154 501840 657160
rect 484216 657076 484268 657082
rect 484216 657018 484268 657024
rect 479524 655716 479576 655722
rect 479524 655658 479576 655664
rect 479536 655602 479564 655658
rect 479536 655574 479826 655602
rect 484228 655588 484256 657018
rect 492956 655852 493008 655858
rect 492956 655794 493008 655800
rect 492968 655588 492996 655794
rect 501800 655588 501828 657154
rect 519358 656024 519414 656033
rect 519358 655959 519414 655968
rect 505836 655648 505888 655654
rect 505888 655596 506230 655602
rect 505836 655590 506230 655596
rect 505848 655574 506230 655590
rect 519372 655588 519400 655959
rect 528112 655588 528140 657455
rect 532514 655888 532570 655897
rect 532514 655823 532570 655832
rect 532528 655588 532556 655823
rect 541360 655588 541388 658310
rect 566464 658300 566516 658306
rect 566464 658242 566516 658248
rect 565176 658232 565228 658238
rect 565176 658174 565228 658180
rect 548616 658164 548668 658170
rect 548616 658106 548668 658112
rect 547142 657248 547198 657257
rect 547142 657183 547198 657192
rect 545764 657008 545816 657014
rect 545764 656950 545816 656956
rect 544476 656600 544528 656606
rect 544476 656542 544528 656548
rect 184848 655444 184900 655450
rect 184848 655386 184900 655392
rect 225328 655376 225380 655382
rect 101982 655314 102180 655330
rect 106398 655314 106688 655330
rect 115230 655314 115520 655330
rect 119554 655314 119936 655330
rect 128386 655314 128768 655330
rect 141542 655314 141832 655330
rect 145958 655314 146248 655330
rect 198568 655314 198674 655330
rect 101982 655308 102192 655314
rect 101982 655302 102140 655308
rect 106398 655308 106700 655314
rect 106398 655302 106648 655308
rect 102140 655250 102192 655256
rect 115230 655308 115532 655314
rect 115230 655302 115480 655308
rect 106648 655250 106700 655256
rect 119554 655308 119948 655314
rect 119554 655302 119896 655308
rect 115480 655250 115532 655256
rect 128386 655308 128780 655314
rect 128386 655302 128728 655308
rect 119896 655250 119948 655256
rect 141542 655308 141844 655314
rect 141542 655302 141792 655308
rect 128728 655250 128780 655256
rect 145958 655308 146260 655314
rect 145958 655302 146208 655308
rect 141792 655250 141844 655256
rect 146208 655250 146260 655256
rect 198556 655308 198674 655314
rect 198608 655302 198674 655308
rect 224986 655324 225328 655330
rect 224986 655318 225380 655324
rect 224986 655302 225368 655318
rect 198556 655250 198608 655256
rect 404820 655240 404872 655246
rect 382936 655178 383226 655194
rect 404872 655188 405122 655194
rect 404820 655182 405122 655188
rect 382924 655172 383226 655178
rect 382976 655166 383226 655172
rect 404832 655166 405122 655182
rect 382924 655114 382976 655120
rect 418160 655104 418212 655110
rect 49514 655072 49570 655081
rect 49266 655030 49514 655058
rect 93490 655072 93546 655081
rect 93242 655030 93490 655058
rect 49514 655007 49570 655016
rect 93490 655007 93546 655016
rect 150254 655072 150310 655081
rect 207570 655072 207626 655081
rect 150310 655030 150374 655058
rect 207414 655030 207570 655058
rect 150254 655007 150310 655016
rect 220910 655072 220966 655081
rect 220662 655030 220910 655058
rect 207570 655007 207626 655016
rect 220910 655007 220966 655016
rect 378506 655072 378562 655081
rect 392122 655072 392178 655081
rect 378562 655030 378810 655058
rect 391966 655030 392122 655058
rect 378506 655007 378562 655016
rect 396092 655042 396382 655058
rect 497002 655072 497058 655081
rect 418212 655052 418370 655058
rect 418160 655046 418370 655052
rect 392122 655007 392178 655016
rect 396080 655036 396382 655042
rect 396132 655030 396382 655036
rect 418172 655030 418370 655046
rect 422496 655042 422694 655058
rect 431144 655042 431526 655058
rect 444392 655042 444682 655058
rect 448808 655042 449098 655058
rect 457456 655042 457838 655058
rect 488552 655042 488658 655058
rect 422484 655036 422694 655042
rect 396080 654978 396132 654984
rect 422536 655030 422694 655036
rect 431132 655036 431526 655042
rect 422484 654978 422536 654984
rect 431184 655030 431526 655036
rect 444380 655036 444682 655042
rect 431132 654978 431184 654984
rect 444432 655030 444682 655036
rect 448796 655036 449098 655042
rect 444380 654978 444432 654984
rect 448848 655030 449098 655036
rect 457444 655036 457838 655042
rect 448796 654978 448848 654984
rect 457496 655030 457838 655036
rect 488540 655036 488658 655042
rect 457444 654978 457496 654984
rect 488592 655030 488658 655036
rect 510250 655072 510306 655081
rect 497058 655030 497398 655058
rect 497002 655007 497058 655016
rect 514758 655072 514814 655081
rect 510306 655030 510554 655058
rect 510250 655007 510306 655016
rect 523590 655072 523646 655081
rect 514814 655030 514970 655058
rect 514758 655007 514814 655016
rect 536838 655072 536894 655081
rect 523646 655030 523802 655058
rect 523590 655007 523646 655016
rect 536894 655030 536958 655058
rect 536838 655007 536894 655016
rect 488540 654978 488592 654984
rect 544384 654560 544436 654566
rect 544384 654502 544436 654508
rect 42248 516112 42300 516118
rect 42248 516054 42300 516060
rect 42156 449880 42208 449886
rect 42156 449822 42208 449828
rect 544396 233238 544424 654502
rect 544488 458182 544516 656542
rect 544476 458176 544528 458182
rect 544476 458118 544528 458124
rect 544384 233232 544436 233238
rect 544384 233174 544436 233180
rect 42064 150408 42116 150414
rect 42064 150350 42116 150356
rect 40684 137964 40736 137970
rect 40684 137906 40736 137912
rect 545776 113150 545804 656950
rect 545856 656736 545908 656742
rect 545856 656678 545908 656684
rect 545868 511970 545896 656678
rect 545856 511964 545908 511970
rect 545856 511906 545908 511912
rect 545764 113144 545816 113150
rect 545764 113086 545816 113092
rect 547156 73166 547184 657183
rect 548524 657144 548576 657150
rect 548524 657086 548576 657092
rect 547236 656804 547288 656810
rect 547236 656746 547288 656752
rect 547248 564398 547276 656746
rect 547236 564392 547288 564398
rect 547236 564334 547288 564340
rect 548536 153202 548564 657086
rect 548628 538218 548656 658106
rect 556896 657960 556948 657966
rect 556896 657902 556948 657908
rect 551376 657892 551428 657898
rect 551376 657834 551428 657840
rect 548708 656872 548760 656878
rect 548708 656814 548760 656820
rect 548720 618254 548748 656814
rect 551282 655616 551338 655625
rect 551282 655551 551338 655560
rect 548708 618248 548760 618254
rect 548708 618190 548760 618196
rect 548616 538212 548668 538218
rect 548616 538154 548668 538160
rect 548524 153196 548576 153202
rect 548524 153138 548576 153144
rect 547144 73160 547196 73166
rect 547144 73102 547196 73108
rect 35808 50108 35860 50114
rect 35808 50050 35860 50056
rect 35164 33108 35216 33114
rect 35164 33050 35216 33056
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 32416 480 32444 3538
rect 33612 480 33640 3538
rect 35820 3398 35848 50050
rect 39948 50040 40000 50046
rect 39948 49982 40000 49988
rect 37188 49292 37240 49298
rect 37188 49234 37240 49240
rect 35992 3732 36044 3738
rect 35992 3674 36044 3680
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 34808 480 34836 3334
rect 36004 480 36032 3674
rect 37200 480 37228 49234
rect 39960 6914 39988 49982
rect 41328 49496 41380 49502
rect 41328 49438 41380 49444
rect 39592 6886 39988 6914
rect 38384 4140 38436 4146
rect 38384 4082 38436 4088
rect 38396 480 38424 4082
rect 39592 480 39620 6886
rect 41340 3398 41368 49438
rect 43272 49230 43300 53108
rect 43444 49904 43496 49910
rect 43444 49846 43496 49852
rect 43260 49224 43312 49230
rect 43260 49166 43312 49172
rect 41880 4072 41932 4078
rect 41880 4014 41932 4020
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 40696 480 40724 3334
rect 41892 480 41920 4014
rect 43456 4010 43484 49846
rect 44284 49366 44312 53108
rect 44824 49836 44876 49842
rect 44824 49778 44876 49784
rect 44272 49360 44324 49366
rect 44272 49302 44324 49308
rect 43444 4004 43496 4010
rect 43444 3946 43496 3952
rect 44836 3806 44864 49778
rect 45296 49026 45324 53108
rect 46308 50386 46336 53108
rect 46296 50380 46348 50386
rect 46296 50322 46348 50328
rect 45468 49972 45520 49978
rect 45468 49914 45520 49920
rect 45284 49020 45336 49026
rect 45284 48962 45336 48968
rect 45376 4004 45428 4010
rect 45376 3946 45428 3952
rect 44824 3800 44876 3806
rect 44824 3742 44876 3748
rect 43076 3664 43128 3670
rect 43076 3606 43128 3612
rect 43088 480 43116 3606
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 44284 480 44312 3334
rect 45388 1986 45416 3946
rect 45480 3398 45508 49914
rect 47320 49774 47348 53108
rect 48332 50454 48360 53108
rect 48320 50448 48372 50454
rect 48320 50390 48372 50396
rect 46204 49768 46256 49774
rect 46204 49710 46256 49716
rect 47308 49768 47360 49774
rect 47308 49710 47360 49716
rect 46216 3466 46244 49710
rect 48228 49224 48280 49230
rect 48228 49166 48280 49172
rect 48240 6914 48268 49166
rect 49344 49094 49372 53108
rect 50356 50522 50384 53108
rect 51368 50726 51396 53108
rect 52380 50862 52408 53108
rect 52472 53094 53406 53122
rect 52368 50856 52420 50862
rect 52368 50798 52420 50804
rect 51356 50720 51408 50726
rect 51356 50662 51408 50668
rect 50344 50516 50396 50522
rect 50344 50458 50396 50464
rect 50988 50448 51040 50454
rect 50988 50390 51040 50396
rect 49608 50380 49660 50386
rect 49608 50322 49660 50328
rect 49332 49088 49384 49094
rect 49332 49030 49384 49036
rect 47872 6886 48268 6914
rect 46664 3800 46716 3806
rect 46664 3742 46716 3748
rect 46204 3460 46256 3466
rect 46204 3402 46256 3408
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45388 1958 45508 1986
rect 45480 480 45508 1958
rect 46676 480 46704 3742
rect 47872 480 47900 6886
rect 49620 3534 49648 50322
rect 50344 49768 50396 49774
rect 50344 49710 50396 49716
rect 50356 4146 50384 49710
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 51000 3534 51028 50390
rect 52368 49360 52420 49366
rect 52368 49302 52420 49308
rect 51080 4548 51132 4554
rect 51080 4490 51132 4496
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51092 3398 51120 4490
rect 52380 3534 52408 49302
rect 52472 4554 52500 53094
rect 54404 50590 54432 53108
rect 54484 50720 54536 50726
rect 54484 50662 54536 50668
rect 54392 50584 54444 50590
rect 54392 50526 54444 50532
rect 53748 50516 53800 50522
rect 53748 50458 53800 50464
rect 52460 4548 52512 4554
rect 52460 4490 52512 4496
rect 53656 4072 53708 4078
rect 53656 4014 53708 4020
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 51080 3392 51132 3398
rect 51080 3334 51132 3340
rect 51368 480 51396 3470
rect 52564 480 52592 3470
rect 53668 2122 53696 4014
rect 53760 3534 53788 50458
rect 54496 3874 54524 50662
rect 55416 50658 55444 53108
rect 56428 50930 56456 53108
rect 56416 50924 56468 50930
rect 56416 50866 56468 50872
rect 57244 50924 57296 50930
rect 57244 50866 57296 50872
rect 56508 50856 56560 50862
rect 56508 50798 56560 50804
rect 55404 50652 55456 50658
rect 55404 50594 55456 50600
rect 55864 50652 55916 50658
rect 55864 50594 55916 50600
rect 55128 49020 55180 49026
rect 55128 48962 55180 48968
rect 55140 6914 55168 48962
rect 54956 6886 55168 6914
rect 54484 3868 54536 3874
rect 54484 3810 54536 3816
rect 53748 3528 53800 3534
rect 53748 3470 53800 3476
rect 53668 2094 53788 2122
rect 53760 480 53788 2094
rect 54956 480 54984 6886
rect 55876 3942 55904 50594
rect 55864 3936 55916 3942
rect 55864 3878 55916 3884
rect 56520 3466 56548 50798
rect 57256 6914 57284 50866
rect 57440 49162 57468 53108
rect 58452 50998 58480 53108
rect 58440 50992 58492 50998
rect 58440 50934 58492 50940
rect 59464 50794 59492 53108
rect 59452 50788 59504 50794
rect 59452 50730 59504 50736
rect 60476 49842 60504 53108
rect 60752 53094 61502 53122
rect 60648 50584 60700 50590
rect 60648 50526 60700 50532
rect 60464 49836 60516 49842
rect 60464 49778 60516 49784
rect 57428 49156 57480 49162
rect 57428 49098 57480 49104
rect 59268 49088 59320 49094
rect 59268 49030 59320 49036
rect 57164 6886 57284 6914
rect 57164 3534 57192 6886
rect 59280 3534 59308 49030
rect 60660 3534 60688 50526
rect 60752 6186 60780 53094
rect 62500 51066 62528 53108
rect 62488 51060 62540 51066
rect 62488 51002 62540 51008
rect 63408 50788 63460 50794
rect 63408 50730 63460 50736
rect 62028 49156 62080 49162
rect 62028 49098 62080 49104
rect 60740 6180 60792 6186
rect 60740 6122 60792 6128
rect 57152 3528 57204 3534
rect 57152 3470 57204 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 60832 3528 60884 3534
rect 60832 3470 60884 3476
rect 56048 3460 56100 3466
rect 56048 3402 56100 3408
rect 56508 3460 56560 3466
rect 56508 3402 56560 3408
rect 56060 480 56088 3402
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57256 480 57284 3266
rect 58452 480 58480 3470
rect 59648 480 59676 3470
rect 60844 480 60872 3470
rect 62040 480 62068 49098
rect 63420 6914 63448 50730
rect 63512 50726 63540 53108
rect 63500 50720 63552 50726
rect 63500 50662 63552 50668
rect 64144 50244 64196 50250
rect 64144 50186 64196 50192
rect 63236 6886 63448 6914
rect 62120 4684 62172 4690
rect 62120 4626 62172 4632
rect 62132 3602 62160 4626
rect 62120 3596 62172 3602
rect 62120 3538 62172 3544
rect 63236 480 63264 6886
rect 64156 4078 64184 50186
rect 64524 50182 64552 53108
rect 64892 53094 65550 53122
rect 64512 50176 64564 50182
rect 64512 50118 64564 50124
rect 64236 49836 64288 49842
rect 64236 49778 64288 49784
rect 64144 4072 64196 4078
rect 64144 4014 64196 4020
rect 64248 3330 64276 49778
rect 64892 4690 64920 53094
rect 66548 50658 66576 53108
rect 67548 50924 67600 50930
rect 67548 50866 67600 50872
rect 66536 50652 66588 50658
rect 66536 50594 66588 50600
rect 66168 49632 66220 49638
rect 66168 49574 66220 49580
rect 64880 4684 64932 4690
rect 64880 4626 64932 4632
rect 64328 3460 64380 3466
rect 64328 3402 64380 3408
rect 64236 3324 64288 3330
rect 64236 3266 64288 3272
rect 64340 480 64368 3402
rect 66180 2922 66208 49574
rect 67560 3602 67588 50866
rect 67652 50862 67680 53108
rect 67744 53094 68678 53122
rect 67640 50856 67692 50862
rect 67640 50798 67692 50804
rect 67744 21418 67772 53094
rect 68928 50856 68980 50862
rect 68928 50798 68980 50804
rect 67732 21412 67784 21418
rect 67732 21354 67784 21360
rect 68940 3602 68968 50798
rect 69676 49910 69704 53108
rect 70308 50924 70360 50930
rect 70308 50866 70360 50872
rect 69664 49904 69716 49910
rect 69664 49846 69716 49852
rect 70216 49564 70268 49570
rect 70216 49506 70268 49512
rect 70228 3602 70256 49506
rect 66720 3596 66772 3602
rect 66720 3538 66772 3544
rect 67548 3596 67600 3602
rect 67548 3538 67600 3544
rect 67916 3596 67968 3602
rect 67916 3538 67968 3544
rect 68928 3596 68980 3602
rect 68928 3538 68980 3544
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 70216 3596 70268 3602
rect 70216 3538 70268 3544
rect 65524 2916 65576 2922
rect 65524 2858 65576 2864
rect 66168 2916 66220 2922
rect 66168 2858 66220 2864
rect 65536 480 65564 2858
rect 66732 480 66760 3538
rect 67928 480 67956 3538
rect 69124 480 69152 3538
rect 70320 480 70348 50866
rect 70688 50318 70716 53108
rect 71044 51060 71096 51066
rect 71044 51002 71096 51008
rect 70676 50312 70728 50318
rect 70676 50254 70728 50260
rect 71056 4010 71084 51002
rect 71136 49904 71188 49910
rect 71136 49846 71188 49852
rect 71044 4004 71096 4010
rect 71044 3946 71096 3952
rect 71148 3738 71176 49846
rect 71700 49434 71728 53108
rect 72712 50114 72740 53108
rect 72700 50108 72752 50114
rect 72700 50050 72752 50056
rect 73724 49910 73752 53108
rect 74448 50244 74500 50250
rect 74448 50186 74500 50192
rect 73712 49904 73764 49910
rect 73712 49846 73764 49852
rect 71688 49428 71740 49434
rect 71688 49370 71740 49376
rect 73068 49428 73120 49434
rect 73068 49370 73120 49376
rect 71504 3936 71556 3942
rect 71504 3878 71556 3884
rect 71136 3732 71188 3738
rect 71136 3674 71188 3680
rect 71516 480 71544 3878
rect 73080 3602 73108 49370
rect 74460 3602 74488 50186
rect 74736 49298 74764 53108
rect 75184 49904 75236 49910
rect 75184 49846 75236 49852
rect 74724 49292 74776 49298
rect 74724 49234 74776 49240
rect 75196 3942 75224 49846
rect 75748 49774 75776 53108
rect 75828 50312 75880 50318
rect 75828 50254 75880 50260
rect 75736 49768 75788 49774
rect 75736 49710 75788 49716
rect 75184 3936 75236 3942
rect 75184 3878 75236 3884
rect 75840 3602 75868 50254
rect 76760 50114 76788 53108
rect 77312 53094 77786 53122
rect 76748 50108 76800 50114
rect 76748 50050 76800 50056
rect 76564 49768 76616 49774
rect 77312 49722 77340 53094
rect 78784 50998 78812 53108
rect 78876 53094 79810 53122
rect 78772 50992 78824 50998
rect 78772 50934 78824 50940
rect 78588 50108 78640 50114
rect 78588 50050 78640 50056
rect 76564 49710 76616 49716
rect 76196 4820 76248 4826
rect 76196 4762 76248 4768
rect 72608 3596 72660 3602
rect 72608 3538 72660 3544
rect 73068 3596 73120 3602
rect 73068 3538 73120 3544
rect 73804 3596 73856 3602
rect 73804 3538 73856 3544
rect 74448 3596 74500 3602
rect 74448 3538 74500 3544
rect 75000 3596 75052 3602
rect 75000 3538 75052 3544
rect 75828 3596 75880 3602
rect 75828 3538 75880 3544
rect 72620 480 72648 3538
rect 73816 480 73844 3538
rect 75012 480 75040 3538
rect 76208 480 76236 4762
rect 76576 3806 76604 49710
rect 77220 49694 77340 49722
rect 77220 49502 77248 49694
rect 77208 49496 77260 49502
rect 77208 49438 77260 49444
rect 76564 3800 76616 3806
rect 76564 3742 76616 3748
rect 78600 3602 78628 50050
rect 78876 3670 78904 53094
rect 80808 49978 80836 53108
rect 81820 51066 81848 53108
rect 81808 51060 81860 51066
rect 81808 51002 81860 51008
rect 81348 50992 81400 50998
rect 81348 50934 81400 50940
rect 80796 49972 80848 49978
rect 80796 49914 80848 49920
rect 79968 49292 80020 49298
rect 79968 49234 80020 49240
rect 79980 6914 80008 49234
rect 79704 6886 80008 6914
rect 78864 3664 78916 3670
rect 78864 3606 78916 3612
rect 77392 3596 77444 3602
rect 77392 3538 77444 3544
rect 78588 3596 78640 3602
rect 78588 3538 78640 3544
rect 77404 480 77432 3538
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 78600 480 78628 3334
rect 79704 480 79732 6886
rect 81360 3602 81388 50934
rect 82084 49972 82136 49978
rect 82084 49914 82136 49920
rect 82096 6914 82124 49914
rect 82832 49774 82860 53108
rect 83464 50040 83516 50046
rect 83464 49982 83516 49988
rect 82820 49768 82872 49774
rect 82820 49710 82872 49716
rect 82004 6886 82124 6914
rect 80888 3596 80940 3602
rect 80888 3538 80940 3544
rect 81348 3596 81400 3602
rect 81348 3538 81400 3544
rect 80900 480 80928 3538
rect 82004 3398 82032 6886
rect 83280 3596 83332 3602
rect 83280 3538 83332 3544
rect 81992 3392 82044 3398
rect 81992 3334 82044 3340
rect 82084 3392 82136 3398
rect 82084 3334 82136 3340
rect 82096 480 82124 3334
rect 83292 480 83320 3538
rect 83476 3398 83504 49982
rect 83844 49230 83872 53108
rect 84856 50386 84884 53108
rect 85868 50454 85896 53108
rect 86512 53094 86894 53122
rect 85856 50448 85908 50454
rect 85856 50390 85908 50396
rect 84844 50380 84896 50386
rect 84844 50322 84896 50328
rect 85488 50108 85540 50114
rect 85488 50050 85540 50056
rect 84108 49496 84160 49502
rect 84108 49438 84160 49444
rect 83832 49224 83884 49230
rect 83832 49166 83884 49172
rect 84120 3602 84148 49438
rect 84108 3596 84160 3602
rect 84108 3538 84160 3544
rect 85500 3534 85528 50050
rect 86512 49366 86540 53094
rect 87892 50522 87920 53108
rect 87880 50516 87932 50522
rect 87880 50458 87932 50464
rect 88248 50380 88300 50386
rect 88248 50322 88300 50328
rect 86868 49836 86920 49842
rect 86868 49778 86920 49784
rect 86500 49360 86552 49366
rect 86500 49302 86552 49308
rect 86776 49224 86828 49230
rect 86776 49166 86828 49172
rect 86788 16574 86816 49166
rect 86696 16546 86816 16574
rect 85672 3596 85724 3602
rect 85672 3538 85724 3544
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 83464 3392 83516 3398
rect 83464 3334 83516 3340
rect 84488 480 84516 3470
rect 85684 480 85712 3538
rect 86696 3482 86724 16546
rect 86880 6914 86908 49778
rect 88260 6914 88288 50322
rect 88904 50182 88932 53108
rect 89076 50720 89128 50726
rect 89076 50662 89128 50668
rect 88892 50176 88944 50182
rect 88892 50118 88944 50124
rect 89088 45554 89116 50662
rect 89916 49026 89944 53108
rect 91020 50590 91048 53108
rect 91008 50584 91060 50590
rect 91008 50526 91060 50532
rect 90364 50448 90416 50454
rect 90364 50390 90416 50396
rect 89904 49020 89956 49026
rect 89904 48962 89956 48968
rect 86788 6886 86908 6914
rect 87984 6886 88288 6914
rect 88996 45526 89116 45554
rect 86788 3602 86816 6886
rect 86776 3596 86828 3602
rect 86776 3538 86828 3544
rect 86696 3454 86908 3482
rect 86880 480 86908 3454
rect 87984 480 88012 6886
rect 88996 3466 89024 45526
rect 90376 6914 90404 50390
rect 92032 49774 92060 53108
rect 92388 50448 92440 50454
rect 92388 50390 92440 50396
rect 92020 49768 92072 49774
rect 92020 49710 92072 49716
rect 91008 49020 91060 49026
rect 91008 48962 91060 48968
rect 90284 6886 90404 6914
rect 90284 3534 90312 6886
rect 91020 3534 91048 48962
rect 92400 3534 92428 50390
rect 93044 49094 93072 53108
rect 94056 50522 94084 53108
rect 95068 50726 95096 53108
rect 95056 50720 95108 50726
rect 95056 50662 95108 50668
rect 95148 50720 95200 50726
rect 95148 50662 95200 50668
rect 94044 50516 94096 50522
rect 94044 50458 94096 50464
rect 93124 49768 93176 49774
rect 93124 49710 93176 49716
rect 93032 49088 93084 49094
rect 93032 49030 93084 49036
rect 92756 4004 92808 4010
rect 92756 3946 92808 3952
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 90272 3528 90324 3534
rect 90272 3470 90324 3476
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 92388 3528 92440 3534
rect 92388 3470 92440 3476
rect 88984 3460 89036 3466
rect 88984 3402 89036 3408
rect 89180 480 89208 3470
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 92768 480 92796 3946
rect 93136 3398 93164 49710
rect 95160 45554 95188 50662
rect 95884 49836 95936 49842
rect 95884 49778 95936 49784
rect 95068 45526 95188 45554
rect 95068 16574 95096 45526
rect 95068 16546 95188 16574
rect 93952 4888 94004 4894
rect 93952 4830 94004 4836
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 93964 480 93992 4830
rect 95160 480 95188 16546
rect 95896 4010 95924 49778
rect 96080 49162 96108 53108
rect 97092 50658 97120 53108
rect 97080 50652 97132 50658
rect 97080 50594 97132 50600
rect 98104 49774 98132 53108
rect 98092 49768 98144 49774
rect 98092 49710 98144 49716
rect 98644 49768 98696 49774
rect 98644 49710 98696 49716
rect 96068 49156 96120 49162
rect 96068 49098 96120 49104
rect 97908 49156 97960 49162
rect 97908 49098 97960 49104
rect 95884 4004 95936 4010
rect 95884 3946 95936 3952
rect 96252 3664 96304 3670
rect 96252 3606 96304 3612
rect 96264 480 96292 3606
rect 97920 3534 97948 49098
rect 98656 3670 98684 49710
rect 99116 49638 99144 53108
rect 100128 50794 100156 53108
rect 101140 50862 101168 53108
rect 101128 50856 101180 50862
rect 101128 50798 101180 50804
rect 100116 50788 100168 50794
rect 100116 50730 100168 50736
rect 99288 50720 99340 50726
rect 99288 50662 99340 50668
rect 99104 49632 99156 49638
rect 99104 49574 99156 49580
rect 98644 3664 98696 3670
rect 98644 3606 98696 3612
rect 99300 3534 99328 50662
rect 100668 50652 100720 50658
rect 100668 50594 100720 50600
rect 100680 3534 100708 50594
rect 102152 49570 102180 53108
rect 103164 50930 103192 53108
rect 103152 50924 103204 50930
rect 103152 50866 103204 50872
rect 103428 50788 103480 50794
rect 103428 50730 103480 50736
rect 102140 49564 102192 49570
rect 102140 49506 102192 49512
rect 102048 49360 102100 49366
rect 102048 49302 102100 49308
rect 102060 3534 102088 49302
rect 103440 3534 103468 50730
rect 104176 49910 104204 53108
rect 104164 49904 104216 49910
rect 104164 49846 104216 49852
rect 105188 49434 105216 53108
rect 106200 50250 106228 53108
rect 107212 50318 107240 53108
rect 107672 53094 108238 53122
rect 107568 50856 107620 50862
rect 107568 50798 107620 50804
rect 107200 50312 107252 50318
rect 107200 50254 107252 50260
rect 106188 50244 106240 50250
rect 106188 50186 106240 50192
rect 106280 50244 106332 50250
rect 106280 50186 106332 50192
rect 106292 50130 106320 50186
rect 106200 50102 106320 50130
rect 105176 49428 105228 49434
rect 105176 49370 105228 49376
rect 104808 49088 104860 49094
rect 104808 49030 104860 49036
rect 104820 6914 104848 49030
rect 104544 6886 104848 6914
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 102232 3528 102284 3534
rect 102232 3470 102284 3476
rect 103428 3528 103480 3534
rect 103428 3470 103480 3476
rect 97460 480 97488 3470
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 101048 480 101076 3470
rect 102244 480 102272 3470
rect 103336 3460 103388 3466
rect 103336 3402 103388 3408
rect 103348 480 103376 3402
rect 104544 480 104572 6886
rect 106200 3534 106228 50102
rect 106924 49904 106976 49910
rect 106924 49846 106976 49852
rect 106936 6914 106964 49846
rect 106844 6886 106964 6914
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 105740 480 105768 3470
rect 106844 3466 106872 6886
rect 107580 3534 107608 50798
rect 107672 4826 107700 53094
rect 109236 50998 109264 53108
rect 109224 50992 109276 50998
rect 109224 50934 109276 50940
rect 110248 49978 110276 53108
rect 110328 50924 110380 50930
rect 110328 50866 110380 50872
rect 110236 49972 110288 49978
rect 110236 49914 110288 49920
rect 108948 22772 109000 22778
rect 108948 22714 109000 22720
rect 107660 4820 107712 4826
rect 107660 4762 107712 4768
rect 108960 3534 108988 22714
rect 110340 3534 110368 50866
rect 111260 49298 111288 53108
rect 112272 51066 112300 53108
rect 112260 51060 112312 51066
rect 112260 51002 112312 51008
rect 113088 50992 113140 50998
rect 113088 50934 113140 50940
rect 111708 50312 111760 50318
rect 111708 50254 111760 50260
rect 111248 49292 111300 49298
rect 111248 49234 111300 49240
rect 111720 3534 111748 50254
rect 113100 6914 113128 50934
rect 113284 50182 113312 53108
rect 113272 50176 113324 50182
rect 113272 50118 113324 50124
rect 114296 49502 114324 53108
rect 115400 50114 115428 53108
rect 115848 51060 115900 51066
rect 115848 51002 115900 51008
rect 115388 50108 115440 50114
rect 115388 50050 115440 50056
rect 114284 49496 114336 49502
rect 114284 49438 114336 49444
rect 112824 6886 113128 6914
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 110328 3528 110380 3534
rect 110328 3470 110380 3476
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 111708 3528 111760 3534
rect 111708 3470 111760 3476
rect 106832 3460 106884 3466
rect 106832 3402 106884 3408
rect 106936 480 106964 3470
rect 108132 480 108160 3470
rect 109328 480 109356 3470
rect 110524 480 110552 3470
rect 111616 3460 111668 3466
rect 111616 3402 111668 3408
rect 111628 480 111656 3402
rect 112824 480 112852 6886
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 114020 480 114048 3538
rect 115860 3534 115888 51002
rect 116412 50046 116440 53108
rect 117228 50176 117280 50182
rect 117228 50118 117280 50124
rect 116400 50040 116452 50046
rect 116400 49982 116452 49988
rect 117240 3534 117268 50118
rect 117424 49230 117452 53108
rect 118436 50522 118464 53108
rect 119448 50590 119476 53108
rect 119436 50584 119488 50590
rect 119436 50526 119488 50532
rect 119988 50584 120040 50590
rect 119988 50526 120040 50532
rect 118424 50516 118476 50522
rect 118424 50458 118476 50464
rect 118608 50108 118660 50114
rect 118608 50050 118660 50056
rect 117412 49224 117464 49230
rect 117412 49166 117464 49172
rect 118620 3534 118648 50050
rect 119896 49972 119948 49978
rect 119896 49914 119948 49920
rect 119908 16574 119936 49914
rect 119816 16546 119936 16574
rect 119816 3534 119844 16546
rect 120000 6914 120028 50526
rect 120460 49026 120488 53108
rect 121368 50516 121420 50522
rect 121368 50458 121420 50464
rect 120448 49020 120500 49026
rect 120448 48962 120500 48968
rect 121380 6914 121408 50458
rect 121472 50454 121500 53108
rect 121460 50448 121512 50454
rect 121460 50390 121512 50396
rect 122484 49842 122512 53108
rect 122852 53094 123510 53122
rect 122748 50448 122800 50454
rect 122748 50390 122800 50396
rect 122472 49836 122524 49842
rect 122472 49778 122524 49784
rect 119908 6886 120028 6914
rect 121104 6886 121408 6914
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 117228 3528 117280 3534
rect 117228 3470 117280 3476
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 118608 3528 118660 3534
rect 118608 3470 118660 3476
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 119804 3528 119856 3534
rect 119804 3470 119856 3476
rect 115216 480 115244 3470
rect 116412 480 116440 3470
rect 117608 480 117636 3470
rect 118804 480 118832 3470
rect 119908 480 119936 6886
rect 121104 480 121132 6886
rect 122760 3330 122788 50390
rect 122852 4894 122880 53094
rect 124508 50386 124536 53108
rect 125152 53094 125534 53122
rect 124496 50380 124548 50386
rect 124496 50322 124548 50328
rect 125152 49910 125180 53094
rect 125508 50040 125560 50046
rect 125508 49982 125560 49988
rect 125140 49904 125192 49910
rect 125140 49846 125192 49852
rect 124128 49836 124180 49842
rect 124128 49778 124180 49784
rect 122840 4888 122892 4894
rect 122840 4830 122892 4836
rect 124140 3534 124168 49778
rect 124864 49768 124916 49774
rect 124864 49710 124916 49716
rect 124876 3602 124904 49710
rect 124864 3596 124916 3602
rect 124864 3538 124916 3544
rect 125520 3534 125548 49982
rect 126532 49162 126560 53108
rect 127544 50726 127572 53108
rect 127532 50720 127584 50726
rect 127532 50662 127584 50668
rect 128556 50658 128584 53108
rect 128544 50652 128596 50658
rect 128544 50594 128596 50600
rect 129568 49366 129596 53108
rect 130580 50794 130608 53108
rect 130568 50788 130620 50794
rect 130568 50730 130620 50736
rect 131592 50386 131620 53108
rect 131580 50380 131632 50386
rect 131580 50322 131632 50328
rect 132408 50380 132460 50386
rect 132408 50322 132460 50328
rect 129556 49360 129608 49366
rect 129556 49302 129608 49308
rect 129004 49292 129056 49298
rect 129004 49234 129056 49240
rect 126520 49156 126572 49162
rect 126520 49098 126572 49104
rect 126888 49020 126940 49026
rect 126888 48962 126940 48968
rect 126900 3534 126928 48962
rect 129016 3534 129044 49234
rect 131028 49224 131080 49230
rect 131028 49166 131080 49172
rect 129648 49156 129700 49162
rect 129648 49098 129700 49104
rect 129660 6914 129688 49098
rect 129384 6886 129688 6914
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 129004 3528 129056 3534
rect 129004 3470 129056 3476
rect 122288 3324 122340 3330
rect 122288 3266 122340 3272
rect 122748 3324 122800 3330
rect 122748 3266 122800 3272
rect 122300 480 122328 3266
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 126992 480 127020 3470
rect 128176 3460 128228 3466
rect 128176 3402 128228 3408
rect 128188 480 128216 3402
rect 129384 480 129412 6886
rect 131040 3534 131068 49166
rect 130568 3528 130620 3534
rect 130568 3470 130620 3476
rect 131028 3528 131080 3534
rect 131028 3470 131080 3476
rect 130580 480 130608 3470
rect 132420 3330 132448 50322
rect 132604 49094 132632 53108
rect 133616 50250 133644 53108
rect 134628 50862 134656 53108
rect 134616 50856 134668 50862
rect 134616 50798 134668 50804
rect 135168 50652 135220 50658
rect 135168 50594 135220 50600
rect 133604 50244 133656 50250
rect 133604 50186 133656 50192
rect 134524 50244 134576 50250
rect 134524 50186 134576 50192
rect 132592 49088 132644 49094
rect 132592 49030 132644 49036
rect 133788 49088 133840 49094
rect 133788 49030 133840 49036
rect 131764 3324 131816 3330
rect 131764 3266 131816 3272
rect 132408 3324 132460 3330
rect 132408 3266 132460 3272
rect 131776 480 131804 3266
rect 133800 3262 133828 49030
rect 134536 22778 134564 50186
rect 134524 22772 134576 22778
rect 134524 22714 134576 22720
rect 135180 3466 135208 50594
rect 135640 50250 135668 53108
rect 136652 50930 136680 53108
rect 136640 50924 136692 50930
rect 136640 50866 136692 50872
rect 136548 50720 136600 50726
rect 136548 50662 136600 50668
rect 135628 50244 135680 50250
rect 135628 50186 135680 50192
rect 136456 3596 136508 3602
rect 136456 3538 136508 3544
rect 134156 3460 134208 3466
rect 134156 3402 134208 3408
rect 135168 3460 135220 3466
rect 135168 3402 135220 3408
rect 132960 3256 133012 3262
rect 132960 3198 133012 3204
rect 133788 3256 133840 3262
rect 133788 3198 133840 3204
rect 132972 480 133000 3198
rect 134168 480 134196 3402
rect 135260 3052 135312 3058
rect 135260 2994 135312 3000
rect 135272 480 135300 2994
rect 136468 480 136496 3538
rect 136560 3058 136588 50662
rect 137664 50318 137692 53108
rect 137928 50788 137980 50794
rect 137928 50730 137980 50736
rect 137652 50312 137704 50318
rect 137652 50254 137704 50260
rect 137284 49768 137336 49774
rect 137284 49710 137336 49716
rect 137296 3398 137324 49710
rect 137940 6914 137968 50730
rect 138768 49774 138796 53108
rect 139780 50998 139808 53108
rect 139768 50992 139820 50998
rect 139768 50934 139820 50940
rect 140688 50992 140740 50998
rect 140688 50934 140740 50940
rect 139308 50924 139360 50930
rect 139308 50866 139360 50872
rect 138756 49768 138808 49774
rect 138756 49710 138808 49716
rect 137664 6886 137968 6914
rect 137284 3392 137336 3398
rect 137284 3334 137336 3340
rect 136548 3052 136600 3058
rect 136548 2994 136600 3000
rect 137664 480 137692 6886
rect 139320 3466 139348 50866
rect 138848 3460 138900 3466
rect 138848 3402 138900 3408
rect 139308 3460 139360 3466
rect 139308 3402 139360 3408
rect 138860 480 138888 3402
rect 140700 3058 140728 50934
rect 140792 49910 140820 53108
rect 141804 51066 141832 53108
rect 141792 51060 141844 51066
rect 141792 51002 141844 51008
rect 142068 50244 142120 50250
rect 142068 50186 142120 50192
rect 140780 49904 140832 49910
rect 140780 49846 140832 49852
rect 142080 3466 142108 50186
rect 142816 50182 142844 53108
rect 143448 50312 143500 50318
rect 143448 50254 143500 50260
rect 142804 50176 142856 50182
rect 142804 50118 142856 50124
rect 143460 3534 143488 50254
rect 143828 50114 143856 53108
rect 144644 51060 144696 51066
rect 144644 51002 144696 51008
rect 143816 50108 143868 50114
rect 143816 50050 143868 50056
rect 144656 45554 144684 51002
rect 144736 50856 144788 50862
rect 144736 50798 144788 50804
rect 144748 48226 144776 50798
rect 144840 49978 144868 53108
rect 145852 50590 145880 53108
rect 145840 50584 145892 50590
rect 145840 50526 145892 50532
rect 146864 50522 146892 53108
rect 146944 50584 146996 50590
rect 146944 50526 146996 50532
rect 146852 50516 146904 50522
rect 146852 50458 146904 50464
rect 144828 49972 144880 49978
rect 144828 49914 144880 49920
rect 146208 49904 146260 49910
rect 146208 49846 146260 49852
rect 144748 48198 144868 48226
rect 144656 45526 144776 45554
rect 144748 16574 144776 45526
rect 144656 16546 144776 16574
rect 144656 3534 144684 16546
rect 144840 6914 144868 48198
rect 146220 6914 146248 49846
rect 144748 6886 144868 6914
rect 145944 6886 146248 6914
rect 142436 3528 142488 3534
rect 142436 3470 142488 3476
rect 143448 3528 143500 3534
rect 143448 3470 143500 3476
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144644 3528 144696 3534
rect 144644 3470 144696 3476
rect 141240 3460 141292 3466
rect 141240 3402 141292 3408
rect 142068 3460 142120 3466
rect 142068 3402 142120 3408
rect 140044 3052 140096 3058
rect 140044 2994 140096 3000
rect 140688 3052 140740 3058
rect 140688 2994 140740 3000
rect 140056 480 140084 2994
rect 141252 480 141280 3402
rect 142448 480 142476 3470
rect 143552 480 143580 3470
rect 144748 480 144776 6886
rect 145944 480 145972 6886
rect 146956 3602 146984 50526
rect 147876 50454 147904 53108
rect 147864 50448 147916 50454
rect 147864 50390 147916 50396
rect 147588 50108 147640 50114
rect 147588 50050 147640 50056
rect 146944 3596 146996 3602
rect 146944 3538 146996 3544
rect 147600 3534 147628 50050
rect 148888 49842 148916 53108
rect 148968 50516 149020 50522
rect 148968 50458 149020 50464
rect 148876 49836 148928 49842
rect 148876 49778 148928 49784
rect 148980 3534 149008 50458
rect 149900 50046 149928 53108
rect 150348 50176 150400 50182
rect 150348 50118 150400 50124
rect 149888 50040 149940 50046
rect 149888 49982 149940 49988
rect 150360 3534 150388 50118
rect 150912 49026 150940 53108
rect 151728 49972 151780 49978
rect 151728 49914 151780 49920
rect 150900 49020 150952 49026
rect 150900 48962 150952 48968
rect 151084 10328 151136 10334
rect 151084 10270 151136 10276
rect 151096 3670 151124 10270
rect 151084 3664 151136 3670
rect 151084 3606 151136 3612
rect 151740 3534 151768 49914
rect 151924 49298 151952 53108
rect 152936 50590 152964 53108
rect 152924 50584 152976 50590
rect 152924 50526 152976 50532
rect 153016 50448 153068 50454
rect 153016 50390 153068 50396
rect 151912 49292 151964 49298
rect 151912 49234 151964 49240
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 150348 3528 150400 3534
rect 150348 3470 150400 3476
rect 150624 3528 150676 3534
rect 150624 3470 150676 3476
rect 151728 3528 151780 3534
rect 151728 3470 151780 3476
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 147140 480 147168 3470
rect 148336 480 148364 3470
rect 149532 480 149560 3470
rect 150636 480 150664 3470
rect 151832 480 151860 3470
rect 153028 480 153056 50390
rect 153108 49904 153160 49910
rect 153108 49846 153160 49852
rect 153120 3534 153148 49846
rect 153948 49162 153976 53108
rect 154488 50040 154540 50046
rect 154488 49982 154540 49988
rect 153936 49156 153988 49162
rect 153936 49098 153988 49104
rect 154500 6914 154528 49982
rect 154960 49230 154988 53108
rect 155972 50386 156000 53108
rect 155960 50380 156012 50386
rect 155960 50322 156012 50328
rect 155868 49836 155920 49842
rect 155868 49778 155920 49784
rect 154948 49224 155000 49230
rect 154948 49166 155000 49172
rect 154224 6886 154528 6914
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 154224 480 154252 6886
rect 155880 3534 155908 49778
rect 156984 49094 157012 53108
rect 157996 50658 158024 53108
rect 159008 50726 159036 53108
rect 159100 53094 160034 53122
rect 158996 50720 159048 50726
rect 158996 50662 159048 50668
rect 157984 50652 158036 50658
rect 157984 50594 158036 50600
rect 158628 50380 158680 50386
rect 158628 50322 158680 50328
rect 157248 49768 157300 49774
rect 157248 49710 157300 49716
rect 156972 49088 157024 49094
rect 156972 49030 157024 49036
rect 157260 3534 157288 49710
rect 158640 3534 158668 50322
rect 159100 45554 159128 53094
rect 161032 50794 161060 53108
rect 162044 50930 162072 53108
rect 163148 50998 163176 53108
rect 163792 53094 164174 53122
rect 163136 50992 163188 50998
rect 163136 50934 163188 50940
rect 162032 50924 162084 50930
rect 162032 50866 162084 50872
rect 161020 50788 161072 50794
rect 161020 50730 161072 50736
rect 161388 50788 161440 50794
rect 161388 50730 161440 50736
rect 160008 50720 160060 50726
rect 160008 50662 160060 50668
rect 158824 45526 159128 45554
rect 158824 10334 158852 45526
rect 158812 10328 158864 10334
rect 158812 10270 158864 10276
rect 160020 3534 160048 50662
rect 161400 3534 161428 50730
rect 162768 50652 162820 50658
rect 162768 50594 162820 50600
rect 162780 6914 162808 50594
rect 163792 50250 163820 53094
rect 165172 50318 165200 53108
rect 166184 51066 166212 53108
rect 166172 51060 166224 51066
rect 166172 51002 166224 51008
rect 165528 50924 165580 50930
rect 165528 50866 165580 50872
rect 165160 50312 165212 50318
rect 165160 50254 165212 50260
rect 163780 50244 163832 50250
rect 163780 50186 163832 50192
rect 164148 50244 164200 50250
rect 164148 50186 164200 50192
rect 162504 6886 162808 6914
rect 155408 3528 155460 3534
rect 155408 3470 155460 3476
rect 155868 3528 155920 3534
rect 155868 3470 155920 3476
rect 156604 3528 156656 3534
rect 156604 3470 156656 3476
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 157800 3528 157852 3534
rect 157800 3470 157852 3476
rect 158628 3528 158680 3534
rect 158628 3470 158680 3476
rect 158904 3528 158956 3534
rect 158904 3470 158956 3476
rect 160008 3528 160060 3534
rect 160008 3470 160060 3476
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 161388 3528 161440 3534
rect 161388 3470 161440 3476
rect 155420 480 155448 3470
rect 156616 480 156644 3470
rect 157812 480 157840 3470
rect 158916 480 158944 3470
rect 160112 480 160140 3470
rect 161296 3460 161348 3466
rect 161296 3402 161348 3408
rect 161308 480 161336 3402
rect 162504 480 162532 6886
rect 164160 3534 164188 50186
rect 163688 3528 163740 3534
rect 163688 3470 163740 3476
rect 164148 3528 164200 3534
rect 164148 3470 164200 3476
rect 163700 480 163728 3470
rect 165540 3058 165568 50866
rect 167196 50862 167224 53108
rect 167184 50856 167236 50862
rect 167184 50798 167236 50804
rect 166908 50720 166960 50726
rect 166908 50662 166960 50668
rect 166920 3534 166948 50662
rect 168208 50590 168236 53108
rect 168288 51060 168340 51066
rect 168288 51002 168340 51008
rect 168196 50584 168248 50590
rect 168196 50526 168248 50532
rect 168300 3534 168328 51002
rect 169220 50114 169248 53108
rect 169668 50584 169720 50590
rect 169668 50526 169720 50532
rect 169576 50312 169628 50318
rect 169576 50254 169628 50260
rect 169208 50108 169260 50114
rect 169208 50050 169260 50056
rect 169588 16574 169616 50254
rect 169496 16546 169616 16574
rect 169496 3534 169524 16546
rect 169680 6914 169708 50526
rect 170232 50522 170260 53108
rect 170220 50516 170272 50522
rect 170220 50458 170272 50464
rect 171048 50516 171100 50522
rect 171048 50458 171100 50464
rect 171060 6914 171088 50458
rect 171244 50182 171272 53108
rect 171232 50176 171284 50182
rect 171232 50118 171284 50124
rect 172256 49978 172284 53108
rect 172244 49972 172296 49978
rect 172244 49914 172296 49920
rect 173268 49910 173296 53108
rect 174280 50454 174308 53108
rect 174268 50448 174320 50454
rect 174268 50390 174320 50396
rect 175188 50176 175240 50182
rect 175188 50118 175240 50124
rect 173808 49972 173860 49978
rect 173808 49914 173860 49920
rect 173256 49904 173308 49910
rect 173256 49846 173308 49852
rect 172428 49768 172480 49774
rect 172428 49710 172480 49716
rect 169588 6886 169708 6914
rect 170784 6886 171088 6914
rect 166080 3528 166132 3534
rect 166080 3470 166132 3476
rect 166908 3528 166960 3534
rect 166908 3470 166960 3476
rect 167184 3528 167236 3534
rect 167184 3470 167236 3476
rect 168288 3528 168340 3534
rect 168288 3470 168340 3476
rect 168380 3528 168432 3534
rect 168380 3470 168432 3476
rect 169484 3528 169536 3534
rect 169484 3470 169536 3476
rect 164884 3052 164936 3058
rect 164884 2994 164936 3000
rect 165528 3052 165580 3058
rect 165528 2994 165580 3000
rect 164896 480 164924 2994
rect 166092 480 166120 3470
rect 167196 480 167224 3470
rect 168392 480 168420 3470
rect 169588 480 169616 6886
rect 170784 480 170812 6886
rect 172440 3534 172468 49710
rect 173820 3534 173848 49914
rect 175200 3534 175228 50118
rect 175292 50046 175320 53108
rect 175280 50040 175332 50046
rect 175280 49982 175332 49988
rect 176304 49842 176332 53108
rect 176568 50108 176620 50114
rect 176568 50050 176620 50056
rect 176292 49836 176344 49842
rect 176292 49778 176344 49784
rect 176580 3534 176608 50050
rect 177316 49910 177344 53108
rect 177856 50448 177908 50454
rect 177856 50390 177908 50396
rect 177304 49904 177356 49910
rect 177304 49846 177356 49852
rect 177868 16574 177896 50390
rect 178328 50386 178356 53108
rect 179340 50862 179368 53108
rect 179328 50856 179380 50862
rect 179328 50798 179380 50804
rect 180064 50856 180116 50862
rect 180064 50798 180116 50804
rect 178316 50380 178368 50386
rect 178316 50322 178368 50328
rect 179328 50380 179380 50386
rect 179328 50322 179380 50328
rect 177948 50040 178000 50046
rect 177948 49982 178000 49988
rect 177776 16546 177896 16574
rect 177776 3534 177804 16546
rect 177960 6914 177988 49982
rect 179340 6914 179368 50322
rect 177868 6886 177988 6914
rect 179064 6886 179368 6914
rect 171968 3528 172020 3534
rect 171968 3470 172020 3476
rect 172428 3528 172480 3534
rect 172428 3470 172480 3476
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 175188 3528 175240 3534
rect 175188 3470 175240 3476
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 176568 3528 176620 3534
rect 176568 3470 176620 3476
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 177764 3528 177816 3534
rect 177764 3470 177816 3476
rect 171980 480 172008 3470
rect 173176 480 173204 3470
rect 174280 480 174308 3470
rect 175476 480 175504 3470
rect 176672 480 176700 3470
rect 177868 480 177896 6886
rect 179064 480 179092 6886
rect 180076 3466 180104 50798
rect 180352 50794 180380 53108
rect 181364 50794 181392 53108
rect 182376 50998 182404 53108
rect 182364 50992 182416 50998
rect 182364 50934 182416 50940
rect 180340 50788 180392 50794
rect 180340 50730 180392 50736
rect 181352 50788 181404 50794
rect 181352 50730 181404 50736
rect 180708 50652 180760 50658
rect 180708 50594 180760 50600
rect 180720 3534 180748 50594
rect 183388 50250 183416 53108
rect 183468 50992 183520 50998
rect 183468 50934 183520 50940
rect 183376 50244 183428 50250
rect 183376 50186 183428 50192
rect 182088 49904 182140 49910
rect 182088 49846 182140 49852
rect 182100 3534 182128 49846
rect 183480 3534 183508 50934
rect 184400 50930 184428 53108
rect 184388 50924 184440 50930
rect 184388 50866 184440 50872
rect 185412 50726 185440 53108
rect 186516 51066 186544 53108
rect 186504 51060 186556 51066
rect 186504 51002 186556 51008
rect 186228 50924 186280 50930
rect 186228 50866 186280 50872
rect 185400 50720 185452 50726
rect 185400 50662 185452 50668
rect 186136 50652 186188 50658
rect 186136 50594 186188 50600
rect 184848 50244 184900 50250
rect 184848 50186 184900 50192
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 181444 3528 181496 3534
rect 181444 3470 181496 3476
rect 182088 3528 182140 3534
rect 182088 3470 182140 3476
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 180064 3460 180116 3466
rect 180064 3402 180116 3408
rect 180260 480 180288 3470
rect 181456 480 181484 3470
rect 182560 480 182588 3470
rect 184860 3262 184888 50186
rect 184940 3528 184992 3534
rect 184940 3470 184992 3476
rect 183744 3256 183796 3262
rect 183744 3198 183796 3204
rect 184848 3256 184900 3262
rect 184848 3198 184900 3204
rect 183756 480 183784 3198
rect 184952 480 184980 3470
rect 186148 480 186176 50594
rect 186240 3534 186268 50866
rect 187528 50318 187556 53108
rect 187608 50720 187660 50726
rect 187608 50662 187660 50668
rect 187516 50312 187568 50318
rect 187516 50254 187568 50260
rect 187620 6914 187648 50662
rect 188540 50590 188568 53108
rect 188528 50584 188580 50590
rect 188528 50526 188580 50532
rect 188988 50584 189040 50590
rect 188988 50526 189040 50532
rect 187344 6886 187648 6914
rect 186228 3528 186280 3534
rect 186228 3470 186280 3476
rect 187344 480 187372 6886
rect 189000 3534 189028 50526
rect 189552 50522 189580 53108
rect 190368 51060 190420 51066
rect 190368 51002 190420 51008
rect 189540 50516 189592 50522
rect 189540 50458 189592 50464
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 188988 3528 189040 3534
rect 188988 3470 189040 3476
rect 188540 480 188568 3470
rect 190380 3466 190408 51002
rect 190564 50862 190592 53108
rect 190552 50856 190604 50862
rect 190552 50798 190604 50804
rect 191576 49978 191604 53108
rect 191748 50312 191800 50318
rect 191748 50254 191800 50260
rect 191564 49972 191616 49978
rect 191564 49914 191616 49920
rect 191760 3534 191788 50254
rect 192588 50182 192616 53108
rect 192576 50176 192628 50182
rect 192576 50118 192628 50124
rect 193600 50114 193628 53108
rect 194416 50856 194468 50862
rect 194416 50798 194468 50804
rect 193588 50108 193640 50114
rect 193588 50050 193640 50056
rect 193128 49972 193180 49978
rect 193128 49914 193180 49920
rect 193140 3534 193168 49914
rect 194428 16574 194456 50798
rect 194508 50516 194560 50522
rect 194508 50458 194560 50464
rect 194336 16546 194456 16574
rect 194336 3534 194364 16546
rect 194520 6914 194548 50458
rect 194612 50454 194640 53108
rect 194600 50448 194652 50454
rect 194600 50390 194652 50396
rect 195624 50046 195652 53108
rect 196636 50386 196664 53108
rect 197648 50794 197676 53108
rect 198384 53094 198674 53122
rect 197636 50788 197688 50794
rect 197636 50730 197688 50736
rect 197268 50448 197320 50454
rect 197268 50390 197320 50396
rect 196624 50380 196676 50386
rect 196624 50322 196676 50328
rect 195888 50176 195940 50182
rect 195888 50118 195940 50124
rect 195612 50040 195664 50046
rect 195612 49982 195664 49988
rect 195900 6914 195928 50118
rect 194428 6886 194548 6914
rect 195624 6886 195928 6914
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 191748 3528 191800 3534
rect 191748 3470 191800 3476
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 193128 3528 193180 3534
rect 193128 3470 193180 3476
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 194324 3528 194376 3534
rect 194324 3470 194376 3476
rect 189724 3460 189776 3466
rect 189724 3402 189776 3408
rect 190368 3460 190420 3466
rect 190368 3402 190420 3408
rect 189736 480 189764 3402
rect 190840 480 190868 3470
rect 192036 480 192064 3470
rect 193232 480 193260 3470
rect 194428 480 194456 6886
rect 195624 480 195652 6886
rect 197280 3330 197308 50390
rect 198384 49910 198412 53094
rect 199672 50998 199700 53108
rect 199660 50992 199712 50998
rect 199660 50934 199712 50940
rect 200028 50992 200080 50998
rect 200028 50934 200080 50940
rect 198648 50788 198700 50794
rect 198648 50730 198700 50736
rect 198372 49904 198424 49910
rect 198372 49846 198424 49852
rect 198660 3534 198688 50730
rect 200040 3534 200068 50934
rect 200684 50250 200712 53108
rect 201696 50930 201724 53108
rect 201684 50924 201736 50930
rect 201684 50866 201736 50872
rect 202708 50658 202736 53108
rect 203720 50726 203748 53108
rect 203708 50720 203760 50726
rect 203708 50662 203760 50668
rect 204168 50720 204220 50726
rect 204168 50662 204220 50668
rect 202696 50652 202748 50658
rect 202696 50594 202748 50600
rect 202788 50652 202840 50658
rect 202788 50594 202840 50600
rect 202800 50504 202828 50594
rect 202708 50476 202828 50504
rect 200672 50244 200724 50250
rect 200672 50186 200724 50192
rect 201408 50244 201460 50250
rect 201408 50186 201460 50192
rect 197912 3528 197964 3534
rect 197912 3470 197964 3476
rect 198648 3528 198700 3534
rect 198648 3470 198700 3476
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 200028 3528 200080 3534
rect 200028 3470 200080 3476
rect 196808 3324 196860 3330
rect 196808 3266 196860 3272
rect 197268 3324 197320 3330
rect 197268 3266 197320 3272
rect 196820 480 196848 3266
rect 197924 480 197952 3470
rect 199120 480 199148 3470
rect 201420 3262 201448 50186
rect 202708 16574 202736 50476
rect 202788 50380 202840 50386
rect 202788 50322 202840 50328
rect 202616 16546 202736 16574
rect 200304 3256 200356 3262
rect 200304 3198 200356 3204
rect 201408 3256 201460 3262
rect 201408 3198 201460 3204
rect 200316 480 200344 3198
rect 202616 3058 202644 16546
rect 202800 6914 202828 50322
rect 204180 6914 204208 50662
rect 204732 50590 204760 53108
rect 205744 51066 205772 53108
rect 205732 51060 205784 51066
rect 205732 51002 205784 51008
rect 205548 50924 205600 50930
rect 205548 50866 205600 50872
rect 204720 50584 204772 50590
rect 204720 50526 204772 50532
rect 202708 6886 202828 6914
rect 203904 6886 204208 6914
rect 201500 3052 201552 3058
rect 201500 2994 201552 3000
rect 202604 3052 202656 3058
rect 202604 2994 202656 3000
rect 201512 480 201540 2994
rect 202708 480 202736 6886
rect 203904 480 203932 6886
rect 205560 3534 205588 50866
rect 206756 50318 206784 53108
rect 206928 50584 206980 50590
rect 206928 50526 206980 50532
rect 206744 50312 206796 50318
rect 206744 50254 206796 50260
rect 206940 3534 206968 50526
rect 207768 49978 207796 53108
rect 208308 51060 208360 51066
rect 208308 51002 208360 51008
rect 207756 49972 207808 49978
rect 207756 49914 207808 49920
rect 208320 3534 208348 51002
rect 208780 50862 208808 53108
rect 208768 50856 208820 50862
rect 208768 50798 208820 50804
rect 209792 50522 209820 53108
rect 209780 50516 209832 50522
rect 209780 50458 209832 50464
rect 209688 50312 209740 50318
rect 209688 50254 209740 50260
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 206192 3528 206244 3534
rect 206192 3470 206244 3476
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 207388 3528 207440 3534
rect 207388 3470 207440 3476
rect 208308 3528 208360 3534
rect 208308 3470 208360 3476
rect 205100 480 205128 3470
rect 206204 480 206232 3470
rect 207400 480 207428 3470
rect 209700 3058 209728 50254
rect 210896 50182 210924 53108
rect 211068 50856 211120 50862
rect 211068 50798 211120 50804
rect 210976 50516 211028 50522
rect 210976 50458 211028 50464
rect 210884 50176 210936 50182
rect 210884 50118 210936 50124
rect 209780 3528 209832 3534
rect 209780 3470 209832 3476
rect 208584 3052 208636 3058
rect 208584 2994 208636 3000
rect 209688 3052 209740 3058
rect 209688 2994 209740 3000
rect 208596 480 208624 2994
rect 209792 480 209820 3470
rect 210988 480 211016 50458
rect 211080 3534 211108 50798
rect 211908 50454 211936 53108
rect 212920 50794 212948 53108
rect 213932 50998 213960 53108
rect 213920 50992 213972 50998
rect 213920 50934 213972 50940
rect 212908 50788 212960 50794
rect 212908 50730 212960 50736
rect 213828 50788 213880 50794
rect 213828 50730 213880 50736
rect 211896 50448 211948 50454
rect 211896 50390 211948 50396
rect 212448 50448 212500 50454
rect 212448 50390 212500 50396
rect 212460 6914 212488 50390
rect 212184 6886 212488 6914
rect 211068 3528 211120 3534
rect 211068 3470 211120 3476
rect 212184 480 212212 6886
rect 213840 3534 213868 50730
rect 214944 50250 214972 53108
rect 215208 50992 215260 50998
rect 215208 50934 215260 50940
rect 214932 50244 214984 50250
rect 214932 50186 214984 50192
rect 215220 3534 215248 50934
rect 215956 50658 215984 53108
rect 215944 50652 215996 50658
rect 215944 50594 215996 50600
rect 216588 50652 216640 50658
rect 216588 50594 216640 50600
rect 216600 3534 216628 50594
rect 216968 50386 216996 53108
rect 217980 50726 218008 53108
rect 218992 50930 219020 53108
rect 218980 50924 219032 50930
rect 218980 50866 219032 50872
rect 219256 50924 219308 50930
rect 219256 50866 219308 50872
rect 217968 50720 218020 50726
rect 217968 50662 218020 50668
rect 216956 50380 217008 50386
rect 216956 50322 217008 50328
rect 217968 50380 218020 50386
rect 217968 50322 218020 50328
rect 217980 3534 218008 50322
rect 219268 16574 219296 50866
rect 219348 50720 219400 50726
rect 219348 50662 219400 50668
rect 219176 16546 219296 16574
rect 219176 3534 219204 16546
rect 219360 6914 219388 50662
rect 220004 50590 220032 53108
rect 221016 51066 221044 53108
rect 221004 51060 221056 51066
rect 221004 51002 221056 51008
rect 219992 50584 220044 50590
rect 219992 50526 220044 50532
rect 220728 50584 220780 50590
rect 220728 50526 220780 50532
rect 220740 6914 220768 50526
rect 222028 50318 222056 53108
rect 222108 51060 222160 51066
rect 222108 51002 222160 51008
rect 222016 50312 222068 50318
rect 222016 50254 222068 50260
rect 219268 6886 219388 6914
rect 220464 6886 220768 6914
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213828 3528 213880 3534
rect 213828 3470 213880 3476
rect 214472 3528 214524 3534
rect 214472 3470 214524 3476
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 216864 3528 216916 3534
rect 216864 3470 216916 3476
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 219164 3528 219216 3534
rect 219164 3470 219216 3476
rect 213380 480 213408 3470
rect 214484 480 214512 3470
rect 215680 480 215708 3470
rect 216876 480 216904 3470
rect 218072 480 218100 3470
rect 219268 480 219296 6886
rect 220464 480 220492 6886
rect 222120 3330 222148 51002
rect 223040 50862 223068 53108
rect 223028 50856 223080 50862
rect 223028 50798 223080 50804
rect 223488 50856 223540 50862
rect 223488 50798 223540 50804
rect 223500 3534 223528 50798
rect 224052 50522 224080 53108
rect 224040 50516 224092 50522
rect 224040 50458 224092 50464
rect 224868 50516 224920 50522
rect 224868 50458 224920 50464
rect 224880 3534 224908 50458
rect 225064 50454 225092 53108
rect 226076 50794 226104 53108
rect 227088 50998 227116 53108
rect 227076 50992 227128 50998
rect 227076 50934 227128 50940
rect 227628 50992 227680 50998
rect 227628 50934 227680 50940
rect 226064 50788 226116 50794
rect 226064 50730 226116 50736
rect 226248 50788 226300 50794
rect 226248 50730 226300 50736
rect 225052 50448 225104 50454
rect 225052 50390 225104 50396
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 221556 3324 221608 3330
rect 221556 3266 221608 3272
rect 222108 3324 222160 3330
rect 222108 3266 222160 3272
rect 221568 480 221596 3266
rect 222764 480 222792 3470
rect 223960 480 223988 3470
rect 226260 3262 226288 50730
rect 227536 50448 227588 50454
rect 227536 50390 227588 50396
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 225144 3256 225196 3262
rect 225144 3198 225196 3204
rect 226248 3256 226300 3262
rect 226248 3198 226300 3204
rect 225156 480 225184 3198
rect 226352 480 226380 3470
rect 227548 480 227576 50390
rect 227640 3534 227668 50934
rect 228100 50658 228128 53108
rect 228088 50652 228140 50658
rect 228088 50594 228140 50600
rect 229008 50652 229060 50658
rect 229008 50594 229060 50600
rect 229020 6914 229048 50594
rect 229112 50386 229140 53108
rect 230124 50930 230152 53108
rect 230112 50924 230164 50930
rect 230112 50866 230164 50872
rect 231136 50726 231164 53108
rect 231124 50720 231176 50726
rect 231124 50662 231176 50668
rect 231768 50720 231820 50726
rect 231768 50662 231820 50668
rect 229100 50380 229152 50386
rect 229100 50322 229152 50328
rect 230388 50380 230440 50386
rect 230388 50322 230440 50328
rect 228744 6886 229048 6914
rect 227628 3528 227680 3534
rect 227628 3470 227680 3476
rect 228744 480 228772 6886
rect 230400 3534 230428 50322
rect 231780 3534 231808 50662
rect 232148 50590 232176 53108
rect 233160 51066 233188 53108
rect 233148 51060 233200 51066
rect 233148 51002 233200 51008
rect 234264 50862 234292 53108
rect 234528 50924 234580 50930
rect 234528 50866 234580 50872
rect 234252 50856 234304 50862
rect 234252 50798 234304 50804
rect 232136 50584 232188 50590
rect 232136 50526 232188 50532
rect 233148 50584 233200 50590
rect 233148 50526 233200 50532
rect 233160 3534 233188 50526
rect 234540 3534 234568 50866
rect 235276 50522 235304 53108
rect 235908 50856 235960 50862
rect 235908 50798 235960 50804
rect 235264 50516 235316 50522
rect 235264 50458 235316 50464
rect 235816 50516 235868 50522
rect 235816 50458 235868 50464
rect 229836 3528 229888 3534
rect 229836 3470 229888 3476
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 229848 480 229876 3470
rect 231044 480 231072 3470
rect 232240 480 232268 3470
rect 233436 480 233464 3470
rect 234632 480 234660 3470
rect 235828 480 235856 50458
rect 235920 3534 235948 50798
rect 236288 50794 236316 53108
rect 237300 50998 237328 53108
rect 237288 50992 237340 50998
rect 237288 50934 237340 50940
rect 236276 50788 236328 50794
rect 236276 50730 236328 50736
rect 237288 50788 237340 50794
rect 237288 50730 237340 50736
rect 237300 6914 237328 50730
rect 238312 50454 238340 53108
rect 239324 50658 239352 53108
rect 239312 50652 239364 50658
rect 239312 50594 239364 50600
rect 240048 50652 240100 50658
rect 240048 50594 240100 50600
rect 238300 50448 238352 50454
rect 238300 50390 238352 50396
rect 238668 50448 238720 50454
rect 238668 50390 238720 50396
rect 237024 6886 237328 6914
rect 235908 3528 235960 3534
rect 235908 3470 235960 3476
rect 237024 480 237052 6886
rect 238680 3534 238708 50390
rect 240060 3534 240088 50594
rect 240336 50386 240364 53108
rect 241348 50726 241376 53108
rect 241428 50992 241480 50998
rect 241428 50934 241480 50940
rect 241336 50720 241388 50726
rect 241336 50662 241388 50668
rect 240324 50380 240376 50386
rect 240324 50322 240376 50328
rect 241440 3534 241468 50934
rect 242360 50590 242388 53108
rect 243372 50930 243400 53108
rect 243360 50924 243412 50930
rect 243360 50866 243412 50872
rect 244384 50862 244412 53108
rect 244372 50856 244424 50862
rect 244372 50798 244424 50804
rect 244188 50720 244240 50726
rect 244188 50662 244240 50668
rect 242348 50584 242400 50590
rect 242348 50526 242400 50532
rect 242808 50584 242860 50590
rect 242808 50526 242860 50532
rect 238116 3528 238168 3534
rect 238116 3470 238168 3476
rect 238668 3528 238720 3534
rect 238668 3470 238720 3476
rect 239312 3528 239364 3534
rect 239312 3470 239364 3476
rect 240048 3528 240100 3534
rect 240048 3470 240100 3476
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 238128 480 238156 3470
rect 239324 480 239352 3470
rect 240520 480 240548 3470
rect 242820 3194 242848 50526
rect 244096 50380 244148 50386
rect 244096 50322 244148 50328
rect 244108 16574 244136 50322
rect 244016 16546 244136 16574
rect 244016 3534 244044 16546
rect 244200 6914 244228 50662
rect 245396 50522 245424 53108
rect 246408 50794 246436 53108
rect 246396 50788 246448 50794
rect 246396 50730 246448 50736
rect 246948 50788 247000 50794
rect 246948 50730 247000 50736
rect 245384 50516 245436 50522
rect 245384 50458 245436 50464
rect 245568 50516 245620 50522
rect 245568 50458 245620 50464
rect 244108 6886 244228 6914
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 244004 3528 244056 3534
rect 244004 3470 244056 3476
rect 241704 3188 241756 3194
rect 241704 3130 241756 3136
rect 242808 3188 242860 3194
rect 242808 3130 242860 3136
rect 241716 480 241744 3130
rect 242912 480 242940 3470
rect 244108 480 244136 6886
rect 245212 598 245424 626
rect 245212 480 245240 598
rect 245396 490 245424 598
rect 245580 490 245608 50458
rect 246960 3126 246988 50730
rect 247420 50454 247448 53108
rect 248432 50658 248460 53108
rect 249444 50998 249472 53108
rect 249432 50992 249484 50998
rect 249432 50934 249484 50940
rect 248420 50652 248472 50658
rect 248420 50594 248472 50600
rect 250456 50590 250484 53108
rect 250444 50584 250496 50590
rect 250444 50526 250496 50532
rect 247408 50448 247460 50454
rect 247408 50390 247460 50396
rect 248328 50448 248380 50454
rect 248328 50390 248380 50396
rect 248340 3534 248368 50390
rect 251468 50386 251496 53108
rect 252376 50992 252428 50998
rect 252376 50934 252428 50940
rect 251456 50380 251508 50386
rect 251456 50322 251508 50328
rect 249708 49836 249760 49842
rect 249708 49778 249760 49784
rect 247592 3528 247644 3534
rect 247592 3470 247644 3476
rect 248328 3528 248380 3534
rect 248328 3470 248380 3476
rect 246396 3120 246448 3126
rect 246396 3062 246448 3068
rect 246948 3120 247000 3126
rect 246948 3062 247000 3068
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245396 462 245608 490
rect 246408 480 246436 3062
rect 247604 480 247632 3470
rect 249720 3058 249748 49778
rect 251088 49768 251140 49774
rect 251088 49710 251140 49716
rect 251100 3534 251128 49710
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 248788 3052 248840 3058
rect 248788 2994 248840 3000
rect 249708 3052 249760 3058
rect 249708 2994 249760 3000
rect 248800 480 248828 2994
rect 249996 480 250024 3470
rect 251192 480 251220 3470
rect 252388 480 252416 50934
rect 252480 50726 252508 53108
rect 252468 50720 252520 50726
rect 252468 50662 252520 50668
rect 253492 50522 253520 53108
rect 253848 50924 253900 50930
rect 253848 50866 253900 50872
rect 253480 50516 253532 50522
rect 253480 50458 253532 50464
rect 252468 50380 252520 50386
rect 252468 50322 252520 50328
rect 252480 3534 252508 50322
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 253492 598 253704 626
rect 253492 480 253520 598
rect 253676 490 253704 598
rect 253860 490 253888 50866
rect 254504 50794 254532 53108
rect 254492 50788 254544 50794
rect 254492 50730 254544 50736
rect 255228 50516 255280 50522
rect 255228 50458 255280 50464
rect 255240 3534 255268 50458
rect 255516 50454 255544 53108
rect 255504 50448 255556 50454
rect 255504 50390 255556 50396
rect 256528 49842 256556 53108
rect 256608 50652 256660 50658
rect 256608 50594 256660 50600
rect 256516 49836 256568 49842
rect 256516 49778 256568 49784
rect 256620 3534 256648 50594
rect 257540 49774 257568 53108
rect 257988 50448 258040 50454
rect 257988 50390 258040 50396
rect 257528 49768 257580 49774
rect 257528 49710 257580 49716
rect 258000 3534 258028 50390
rect 258644 50386 258672 53108
rect 259656 50998 259684 53108
rect 259644 50992 259696 50998
rect 259644 50934 259696 50940
rect 260668 50930 260696 53108
rect 260656 50924 260708 50930
rect 260656 50866 260708 50872
rect 261680 50522 261708 53108
rect 262128 50856 262180 50862
rect 262128 50798 262180 50804
rect 261668 50516 261720 50522
rect 261668 50458 261720 50464
rect 258632 50380 258684 50386
rect 258632 50322 258684 50328
rect 260656 49904 260708 49910
rect 260656 49846 260708 49852
rect 259368 49836 259420 49842
rect 259368 49778 259420 49784
rect 259380 3534 259408 49778
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 255228 3528 255280 3534
rect 255228 3470 255280 3476
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 256608 3528 256660 3534
rect 256608 3470 256660 3476
rect 257068 3528 257120 3534
rect 257068 3470 257120 3476
rect 257988 3528 258040 3534
rect 257988 3470 258040 3476
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 253676 462 253888 490
rect 254688 480 254716 3470
rect 255884 480 255912 3470
rect 257080 480 257108 3470
rect 258276 480 258304 3470
rect 259472 480 259500 3470
rect 260668 480 260696 49846
rect 260748 49768 260800 49774
rect 260748 49710 260800 49716
rect 260760 3534 260788 49710
rect 260748 3528 260800 3534
rect 260748 3470 260800 3476
rect 261772 598 261984 626
rect 261772 480 261800 598
rect 261956 490 261984 598
rect 262140 490 262168 50798
rect 262692 50658 262720 53108
rect 262680 50652 262732 50658
rect 262680 50594 262732 50600
rect 263704 50454 263732 53108
rect 263692 50448 263744 50454
rect 263692 50390 263744 50396
rect 263508 50040 263560 50046
rect 263508 49982 263560 49988
rect 263520 3534 263548 49982
rect 264716 49842 264744 53108
rect 264888 50788 264940 50794
rect 264888 50730 264940 50736
rect 264704 49836 264756 49842
rect 264704 49778 264756 49784
rect 264900 3534 264928 50730
rect 265728 49774 265756 53108
rect 266740 49910 266768 53108
rect 267752 50862 267780 53108
rect 267740 50856 267792 50862
rect 267740 50798 267792 50804
rect 267648 50720 267700 50726
rect 267648 50662 267700 50668
rect 267004 50584 267056 50590
rect 267004 50526 267056 50532
rect 266728 49904 266780 49910
rect 266728 49846 266780 49852
rect 265716 49768 265768 49774
rect 265716 49710 265768 49716
rect 262956 3528 263008 3534
rect 262956 3470 263008 3476
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 264888 3528 264940 3534
rect 264888 3470 264940 3476
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 261956 462 262168 490
rect 262968 480 262996 3470
rect 264164 480 264192 3470
rect 265348 3460 265400 3466
rect 265348 3402 265400 3408
rect 265360 480 265388 3402
rect 266556 480 266584 3470
rect 267016 3466 267044 50526
rect 267660 3534 267688 50662
rect 268764 50046 268792 53108
rect 269776 50794 269804 53108
rect 269764 50788 269816 50794
rect 269764 50730 269816 50736
rect 270788 50590 270816 53108
rect 271800 50726 271828 53108
rect 271788 50720 271840 50726
rect 271788 50662 271840 50668
rect 270776 50584 270828 50590
rect 270776 50526 270828 50532
rect 268752 50040 268804 50046
rect 268752 49982 268804 49988
rect 270408 49972 270460 49978
rect 270408 49914 270460 49920
rect 269028 49904 269080 49910
rect 269028 49846 269080 49852
rect 268936 49768 268988 49774
rect 268936 49710 268988 49716
rect 268948 3602 268976 49710
rect 267740 3596 267792 3602
rect 267740 3538 267792 3544
rect 268936 3596 268988 3602
rect 268936 3538 268988 3544
rect 267648 3528 267700 3534
rect 267648 3470 267700 3476
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 267752 480 267780 3538
rect 269040 3482 269068 49846
rect 268856 3454 269068 3482
rect 268856 480 268884 3454
rect 270052 598 270264 626
rect 270052 480 270080 598
rect 270236 490 270264 598
rect 270420 490 270448 49914
rect 271788 49836 271840 49842
rect 271788 49778 271840 49784
rect 271800 3330 271828 49778
rect 272812 49774 272840 53108
rect 273824 49910 273852 53108
rect 274548 50652 274600 50658
rect 274548 50594 274600 50600
rect 273812 49904 273864 49910
rect 273812 49846 273864 49852
rect 272800 49768 272852 49774
rect 272800 49710 272852 49716
rect 273904 49768 273956 49774
rect 273904 49710 273956 49716
rect 273628 3528 273680 3534
rect 273628 3470 273680 3476
rect 272432 3460 272484 3466
rect 272432 3402 272484 3408
rect 271236 3324 271288 3330
rect 271236 3266 271288 3272
rect 271788 3324 271840 3330
rect 271788 3266 271840 3272
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270236 462 270448 490
rect 271248 480 271276 3266
rect 272444 480 272472 3402
rect 273640 480 273668 3470
rect 273916 3466 273944 49710
rect 274560 3534 274588 50594
rect 274836 49978 274864 53108
rect 274824 49972 274876 49978
rect 274824 49914 274876 49920
rect 275848 49842 275876 53108
rect 275928 50788 275980 50794
rect 275928 50730 275980 50736
rect 275836 49836 275888 49842
rect 275836 49778 275888 49784
rect 275940 3534 275968 50730
rect 276860 49774 276888 53108
rect 277308 50720 277360 50726
rect 277308 50662 277360 50668
rect 277216 50380 277268 50386
rect 277216 50322 277268 50328
rect 276848 49768 276900 49774
rect 276848 49710 276900 49716
rect 277228 6914 277256 50322
rect 277136 6886 277256 6914
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 274824 3528 274876 3534
rect 274824 3470 274876 3476
rect 275928 3528 275980 3534
rect 275928 3470 275980 3476
rect 273904 3460 273956 3466
rect 273904 3402 273956 3408
rect 274836 480 274864 3470
rect 276020 3324 276072 3330
rect 276020 3266 276072 3272
rect 276032 480 276060 3266
rect 277136 480 277164 6886
rect 277320 3330 277348 50662
rect 277872 50658 277900 53108
rect 278884 50794 278912 53108
rect 278872 50788 278924 50794
rect 278872 50730 278924 50736
rect 279896 50726 279924 53108
rect 279884 50720 279936 50726
rect 279884 50662 279936 50668
rect 277860 50652 277912 50658
rect 277860 50594 277912 50600
rect 280908 50386 280936 53108
rect 280896 50380 280948 50386
rect 280896 50322 280948 50328
rect 280068 49904 280120 49910
rect 280068 49846 280120 49852
rect 278688 49768 278740 49774
rect 278688 49710 278740 49716
rect 277308 3324 277360 3330
rect 277308 3266 277360 3272
rect 278332 598 278544 626
rect 278332 480 278360 598
rect 278516 490 278544 598
rect 278700 490 278728 49710
rect 280080 3330 280108 49846
rect 281448 49836 281500 49842
rect 281448 49778 281500 49784
rect 281460 3534 281488 49778
rect 282012 49774 282040 53108
rect 283024 49910 283052 53108
rect 283012 49904 283064 49910
rect 283012 49846 283064 49852
rect 284036 49842 284064 53108
rect 284024 49836 284076 49842
rect 284024 49778 284076 49784
rect 285048 49774 285076 53108
rect 285784 53094 286074 53122
rect 285496 50788 285548 50794
rect 285496 50730 285548 50736
rect 282000 49768 282052 49774
rect 282000 49710 282052 49716
rect 282828 49768 282880 49774
rect 282828 49710 282880 49716
rect 285036 49768 285088 49774
rect 285036 49710 285088 49716
rect 282840 3534 282868 49710
rect 285508 6914 285536 50730
rect 285588 50720 285640 50726
rect 285588 50662 285640 50668
rect 285416 6886 285536 6914
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 281908 3528 281960 3534
rect 281908 3470 281960 3476
rect 282828 3528 282880 3534
rect 282828 3470 282880 3476
rect 284300 3528 284352 3534
rect 284300 3470 284352 3476
rect 279516 3324 279568 3330
rect 279516 3266 279568 3272
rect 280068 3324 280120 3330
rect 280068 3266 280120 3272
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 278516 462 278728 490
rect 279528 480 279556 3266
rect 280724 480 280752 3470
rect 281920 480 281948 3470
rect 283104 3188 283156 3194
rect 283104 3130 283156 3136
rect 283116 480 283144 3130
rect 284312 480 284340 3470
rect 285416 480 285444 6886
rect 285600 3534 285628 50662
rect 285588 3528 285640 3534
rect 285588 3470 285640 3476
rect 285784 3194 285812 53094
rect 287072 50726 287100 53108
rect 288084 50794 288112 53108
rect 288072 50788 288124 50794
rect 288072 50730 288124 50736
rect 287060 50720 287112 50726
rect 287060 50662 287112 50668
rect 289096 50590 289124 53108
rect 286968 50584 287020 50590
rect 286968 50526 287020 50532
rect 289084 50584 289136 50590
rect 289084 50526 289136 50532
rect 285772 3188 285824 3194
rect 285772 3130 285824 3136
rect 286612 598 286824 626
rect 286612 480 286640 598
rect 286796 490 286824 598
rect 286980 490 287008 50526
rect 290108 49842 290136 53108
rect 288348 49836 288400 49842
rect 288348 49778 288400 49784
rect 290096 49836 290148 49842
rect 290096 49778 290148 49784
rect 288360 3534 288388 49778
rect 291120 49774 291148 53108
rect 291304 53094 292146 53122
rect 292592 53094 293158 53122
rect 294064 53094 294170 53122
rect 294800 53094 295182 53122
rect 295444 53094 296194 53122
rect 296732 53094 297206 53122
rect 289728 49768 289780 49774
rect 289728 49710 289780 49716
rect 291108 49768 291160 49774
rect 291108 49710 291160 49716
rect 289740 3534 289768 49710
rect 291304 3534 291332 53094
rect 292592 49722 292620 53094
rect 292500 49694 292620 49722
rect 292500 3534 292528 49694
rect 293960 46164 294012 46170
rect 293960 46106 294012 46112
rect 287796 3528 287848 3534
rect 287796 3470 287848 3476
rect 288348 3528 288400 3534
rect 288348 3470 288400 3476
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 291292 3528 291344 3534
rect 291292 3470 291344 3476
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 292488 3528 292540 3534
rect 292488 3470 292540 3476
rect 292580 3528 292632 3534
rect 292580 3470 292632 3476
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 286796 462 287008 490
rect 287808 480 287836 3470
rect 289004 480 289032 3470
rect 290200 480 290228 3470
rect 291396 480 291424 3470
rect 292592 480 292620 3470
rect 293972 2802 294000 46106
rect 294064 3534 294092 53094
rect 294800 46170 294828 53094
rect 294788 46164 294840 46170
rect 294788 46106 294840 46112
rect 294052 3528 294104 3534
rect 294052 3470 294104 3476
rect 295444 2854 295472 53094
rect 296732 50674 296760 53094
rect 296640 50646 296760 50674
rect 296640 3534 296668 50646
rect 298100 49360 298152 49366
rect 298100 49302 298152 49308
rect 296076 3528 296128 3534
rect 296076 3470 296128 3476
rect 296628 3528 296680 3534
rect 296628 3470 296680 3476
rect 293696 2774 294000 2802
rect 294880 2848 294932 2854
rect 294880 2790 294932 2796
rect 295432 2848 295484 2854
rect 295432 2790 295484 2796
rect 293696 480 293724 2774
rect 294892 480 294920 2790
rect 296088 480 296116 3470
rect 297272 3120 297324 3126
rect 297272 3062 297324 3068
rect 297284 480 297312 3062
rect 298112 490 298140 49302
rect 298204 3126 298232 53108
rect 298848 53094 299230 53122
rect 299492 53094 300242 53122
rect 300872 53094 301254 53122
rect 302266 53094 302372 53122
rect 298848 49366 298876 53094
rect 298836 49360 298888 49366
rect 298836 49302 298888 49308
rect 299492 16574 299520 53094
rect 300872 49722 300900 53094
rect 300780 49694 300900 49722
rect 299492 16546 299704 16574
rect 298192 3120 298244 3126
rect 298192 3062 298244 3068
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 16546
rect 300780 480 300808 49694
rect 302344 6914 302372 53094
rect 302252 6886 302372 6914
rect 302436 53094 303278 53122
rect 303632 53094 304290 53122
rect 305012 53094 305302 53122
rect 302252 3482 302280 6886
rect 302436 3534 302464 53094
rect 303632 16574 303660 53094
rect 303632 16546 303936 16574
rect 301976 3454 302280 3482
rect 302424 3528 302476 3534
rect 302424 3470 302476 3476
rect 303160 3528 303212 3534
rect 303160 3470 303212 3476
rect 301976 480 302004 3454
rect 303172 480 303200 3470
rect 303908 490 303936 16546
rect 305012 3330 305040 53094
rect 305000 3324 305052 3330
rect 305000 3266 305052 3272
rect 305552 3324 305604 3330
rect 305552 3266 305604 3272
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3266
rect 306392 490 306420 53108
rect 307418 53094 307708 53122
rect 307680 3346 307708 53094
rect 307772 53094 308430 53122
rect 309152 53094 309442 53122
rect 307772 3534 307800 53094
rect 307760 3528 307812 3534
rect 307760 3470 307812 3476
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 307680 3318 307984 3346
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 3318
rect 309060 480 309088 3470
rect 309152 3262 309180 53094
rect 310440 3534 310468 53108
rect 311466 53094 311848 53122
rect 311820 3534 311848 53094
rect 312464 49774 312492 53108
rect 313476 49910 313504 53108
rect 314502 53094 314608 53122
rect 315514 53094 315896 53122
rect 313464 49904 313516 49910
rect 313464 49846 313516 49852
rect 314476 49904 314528 49910
rect 314476 49846 314528 49852
rect 312452 49768 312504 49774
rect 312452 49710 312504 49716
rect 313464 49768 313516 49774
rect 313464 49710 313516 49716
rect 313476 16574 313504 49710
rect 313476 16546 313872 16574
rect 310428 3528 310480 3534
rect 310428 3470 310480 3476
rect 311440 3528 311492 3534
rect 311440 3470 311492 3476
rect 311808 3528 311860 3534
rect 311808 3470 311860 3476
rect 312636 3528 312688 3534
rect 312636 3470 312688 3476
rect 309140 3256 309192 3262
rect 309140 3198 309192 3204
rect 310244 3256 310296 3262
rect 310244 3198 310296 3204
rect 310256 480 310284 3198
rect 311452 480 311480 3470
rect 312648 480 312676 3470
rect 313844 480 313872 16546
rect 314488 3534 314516 49846
rect 314580 4078 314608 53094
rect 315868 50674 315896 53094
rect 315868 50646 316172 50674
rect 316144 45554 316172 50646
rect 316512 49774 316540 53108
rect 317524 49842 317552 53108
rect 318550 53094 318656 53122
rect 317512 49836 317564 49842
rect 317512 49778 317564 49784
rect 316500 49768 316552 49774
rect 316500 49710 316552 49716
rect 317604 49768 317656 49774
rect 317604 49710 317656 49716
rect 316144 45526 316264 45554
rect 316236 16574 316264 45526
rect 317616 16574 317644 49710
rect 316236 16546 317368 16574
rect 317616 16546 318104 16574
rect 314568 4072 314620 4078
rect 314568 4014 314620 4020
rect 316224 4072 316276 4078
rect 316224 4014 316276 4020
rect 314476 3528 314528 3534
rect 314476 3470 314528 3476
rect 315028 3528 315080 3534
rect 315028 3470 315080 3476
rect 315040 480 315068 3470
rect 316236 480 316264 4014
rect 317340 480 317368 16546
rect 318076 490 318104 16546
rect 318628 3058 318656 53094
rect 319548 49842 319576 53108
rect 318708 49836 318760 49842
rect 318708 49778 318760 49784
rect 319536 49836 319588 49842
rect 319536 49778 319588 49784
rect 318720 3534 318748 49778
rect 320560 49774 320588 53108
rect 320824 49836 320876 49842
rect 320824 49778 320876 49784
rect 320548 49768 320600 49774
rect 320548 49710 320600 49716
rect 318708 3528 318760 3534
rect 318708 3470 318760 3476
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 318616 3052 318668 3058
rect 318616 2994 318668 3000
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 3470
rect 320836 2990 320864 49778
rect 321572 49774 321600 53108
rect 322598 53094 322888 53122
rect 323610 53094 324268 53122
rect 321468 49768 321520 49774
rect 321468 49710 321520 49716
rect 321560 49768 321612 49774
rect 321560 49710 321612 49716
rect 322756 49768 322808 49774
rect 322756 49710 322808 49716
rect 321480 3466 321508 49710
rect 322768 3534 322796 49710
rect 322756 3528 322808 3534
rect 322756 3470 322808 3476
rect 321468 3460 321520 3466
rect 321468 3402 321520 3408
rect 322860 3262 322888 53094
rect 324240 3602 324268 53094
rect 324608 49774 324636 53108
rect 324596 49768 324648 49774
rect 324596 49710 324648 49716
rect 325516 49768 325568 49774
rect 325516 49710 325568 49716
rect 324228 3596 324280 3602
rect 324228 3538 324280 3544
rect 324412 3528 324464 3534
rect 324412 3470 324464 3476
rect 323308 3460 323360 3466
rect 323308 3402 323360 3408
rect 322848 3256 322900 3262
rect 322848 3198 322900 3204
rect 320916 3052 320968 3058
rect 320916 2994 320968 3000
rect 320824 2984 320876 2990
rect 320824 2926 320876 2932
rect 320928 480 320956 2994
rect 322112 2984 322164 2990
rect 322112 2926 322164 2932
rect 322124 480 322152 2926
rect 323320 480 323348 3402
rect 324424 480 324452 3470
rect 325528 3330 325556 49710
rect 325620 3466 325648 53108
rect 326646 53094 327028 53122
rect 327658 53094 328408 53122
rect 326804 3596 326856 3602
rect 326804 3538 326856 3544
rect 325608 3460 325660 3466
rect 325608 3402 325660 3408
rect 325516 3324 325568 3330
rect 325516 3266 325568 3272
rect 325608 3256 325660 3262
rect 325608 3198 325660 3204
rect 325620 480 325648 3198
rect 326816 480 326844 3538
rect 327000 3194 327028 53094
rect 328380 3602 328408 53094
rect 328656 49774 328684 53108
rect 329668 53094 329774 53122
rect 330786 53094 331168 53122
rect 328644 49768 328696 49774
rect 328644 49710 328696 49716
rect 328368 3596 328420 3602
rect 328368 3538 328420 3544
rect 329196 3460 329248 3466
rect 329196 3402 329248 3408
rect 328000 3324 328052 3330
rect 328000 3266 328052 3272
rect 326988 3188 327040 3194
rect 326988 3130 327040 3136
rect 328012 480 328040 3266
rect 329208 480 329236 3402
rect 329668 3398 329696 53094
rect 329748 49768 329800 49774
rect 329748 49710 329800 49716
rect 329760 3534 329788 49710
rect 329748 3528 329800 3534
rect 329748 3470 329800 3476
rect 331140 3466 331168 53094
rect 331784 49774 331812 53108
rect 332796 50794 332824 53108
rect 332784 50788 332836 50794
rect 332784 50730 332836 50736
rect 333808 49774 333836 53108
rect 334834 53094 335308 53122
rect 331772 49768 331824 49774
rect 331772 49710 331824 49716
rect 332508 49768 332560 49774
rect 332508 49710 332560 49716
rect 333796 49768 333848 49774
rect 333796 49710 333848 49716
rect 334624 49768 334676 49774
rect 334624 49710 334676 49716
rect 332520 4078 332548 49710
rect 332508 4072 332560 4078
rect 332508 4014 332560 4020
rect 334636 3602 334664 49710
rect 331588 3596 331640 3602
rect 331588 3538 331640 3544
rect 334624 3596 334676 3602
rect 334624 3538 334676 3544
rect 331128 3460 331180 3466
rect 331128 3402 331180 3408
rect 329656 3392 329708 3398
rect 329656 3334 329708 3340
rect 330392 3188 330444 3194
rect 330392 3130 330444 3136
rect 330404 480 330432 3130
rect 331600 480 331628 3538
rect 335280 3534 335308 53094
rect 335832 49774 335860 53108
rect 336004 50788 336056 50794
rect 336004 50730 336056 50736
rect 335820 49768 335872 49774
rect 335820 49710 335872 49716
rect 336016 3534 336044 50730
rect 336844 49842 336872 53108
rect 336832 49836 336884 49842
rect 336832 49778 336884 49784
rect 337856 49774 337884 53108
rect 338882 53094 339448 53122
rect 338856 49836 338908 49842
rect 338856 49778 338908 49784
rect 336648 49768 336700 49774
rect 336648 49710 336700 49716
rect 337844 49768 337896 49774
rect 337844 49710 337896 49716
rect 338764 49768 338816 49774
rect 338764 49710 338816 49716
rect 336280 4072 336332 4078
rect 336280 4014 336332 4020
rect 332692 3528 332744 3534
rect 332692 3470 332744 3476
rect 335268 3528 335320 3534
rect 335268 3470 335320 3476
rect 336004 3528 336056 3534
rect 336004 3470 336056 3476
rect 332704 480 332732 3470
rect 335084 3460 335136 3466
rect 335084 3402 335136 3408
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 335096 480 335124 3402
rect 336292 480 336320 4014
rect 336660 3262 336688 49710
rect 338672 3596 338724 3602
rect 338672 3538 338724 3544
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 336648 3256 336700 3262
rect 336648 3198 336700 3204
rect 337488 480 337516 3470
rect 338684 480 338712 3538
rect 338776 3534 338804 49710
rect 338764 3528 338816 3534
rect 338764 3470 338816 3476
rect 338868 3330 338896 49778
rect 339420 3602 339448 53094
rect 339880 49774 339908 53108
rect 340892 49774 340920 53108
rect 341918 53094 342116 53122
rect 342930 53094 343588 53122
rect 339868 49768 339920 49774
rect 339868 49710 339920 49716
rect 340788 49768 340840 49774
rect 340788 49710 340840 49716
rect 340880 49768 340932 49774
rect 340880 49710 340932 49716
rect 340800 4078 340828 49710
rect 340788 4072 340840 4078
rect 340788 4014 340840 4020
rect 339408 3596 339460 3602
rect 339408 3538 339460 3544
rect 342088 3466 342116 53094
rect 342168 49768 342220 49774
rect 342168 49710 342220 49716
rect 342180 4146 342208 49710
rect 342168 4140 342220 4146
rect 342168 4082 342220 4088
rect 343560 3670 343588 53094
rect 343928 50386 343956 53108
rect 343916 50380 343968 50386
rect 343916 50322 343968 50328
rect 344940 3806 344968 53108
rect 345966 53094 346348 53122
rect 346978 53094 347728 53122
rect 345756 4072 345808 4078
rect 345756 4014 345808 4020
rect 344928 3800 344980 3806
rect 344928 3742 344980 3748
rect 343548 3664 343600 3670
rect 343548 3606 343600 3612
rect 344560 3596 344612 3602
rect 344560 3538 344612 3544
rect 343364 3528 343416 3534
rect 343364 3470 343416 3476
rect 339868 3460 339920 3466
rect 339868 3402 339920 3408
rect 342076 3460 342128 3466
rect 342076 3402 342128 3408
rect 338856 3324 338908 3330
rect 338856 3266 338908 3272
rect 339880 480 339908 3402
rect 342168 3324 342220 3330
rect 342168 3266 342220 3272
rect 340972 3256 341024 3262
rect 340972 3198 341024 3204
rect 340984 480 341012 3198
rect 342180 480 342208 3266
rect 343376 480 343404 3470
rect 344572 480 344600 3538
rect 345768 480 345796 4014
rect 346320 3058 346348 53094
rect 346952 4140 347004 4146
rect 346952 4082 347004 4088
rect 346308 3052 346360 3058
rect 346308 2994 346360 3000
rect 346964 480 346992 4082
rect 347700 3534 347728 53094
rect 347976 49774 348004 53108
rect 349002 53094 349108 53122
rect 350014 53094 350488 53122
rect 347964 49768 348016 49774
rect 347964 49710 348016 49716
rect 348976 49768 349028 49774
rect 348976 49710 349028 49716
rect 348988 4146 349016 49710
rect 348976 4140 349028 4146
rect 348976 4082 349028 4088
rect 347688 3528 347740 3534
rect 347688 3470 347740 3476
rect 348056 3460 348108 3466
rect 348056 3402 348108 3408
rect 348068 480 348096 3402
rect 349080 2990 349108 53094
rect 349252 50380 349304 50386
rect 349252 50322 349304 50328
rect 349264 16574 349292 50322
rect 349264 16546 350396 16574
rect 349252 3664 349304 3670
rect 349252 3606 349304 3612
rect 349068 2984 349120 2990
rect 349068 2926 349120 2932
rect 349264 480 349292 3606
rect 350368 3482 350396 16546
rect 350460 3738 350488 53094
rect 351012 49774 351040 53108
rect 352024 49774 352052 53108
rect 353050 53094 353248 53122
rect 354154 53094 354628 53122
rect 351000 49768 351052 49774
rect 351000 49710 351052 49716
rect 351828 49768 351880 49774
rect 351828 49710 351880 49716
rect 352012 49768 352064 49774
rect 352012 49710 352064 49716
rect 353116 49768 353168 49774
rect 353116 49710 353168 49716
rect 351840 4078 351868 49710
rect 351828 4072 351880 4078
rect 351828 4014 351880 4020
rect 353128 3874 353156 49710
rect 353220 3942 353248 53094
rect 353208 3936 353260 3942
rect 353208 3878 353260 3884
rect 353116 3868 353168 3874
rect 353116 3810 353168 3816
rect 351644 3800 351696 3806
rect 351644 3742 351696 3748
rect 350448 3732 350500 3738
rect 350448 3674 350500 3680
rect 350368 3454 350488 3482
rect 350460 480 350488 3454
rect 351656 480 351684 3742
rect 354600 3602 354628 53094
rect 355152 49774 355180 53108
rect 356164 49774 356192 53108
rect 357190 53094 357296 53122
rect 358202 53094 358768 53122
rect 355140 49768 355192 49774
rect 355140 49710 355192 49716
rect 355968 49768 356020 49774
rect 355968 49710 356020 49716
rect 356152 49768 356204 49774
rect 356152 49710 356204 49716
rect 355232 4140 355284 4146
rect 355232 4082 355284 4088
rect 354588 3596 354640 3602
rect 354588 3538 354640 3544
rect 354036 3528 354088 3534
rect 354036 3470 354088 3476
rect 352840 3052 352892 3058
rect 352840 2994 352892 3000
rect 352852 480 352880 2994
rect 354048 480 354076 3470
rect 355244 480 355272 4082
rect 355980 3534 356008 49710
rect 357268 3670 357296 53094
rect 357348 49768 357400 49774
rect 357348 49710 357400 49716
rect 357360 4010 357388 49710
rect 358740 6914 358768 53094
rect 359200 49774 359228 53108
rect 360212 49774 360240 53108
rect 361238 53094 361436 53122
rect 362250 53094 362908 53122
rect 359188 49768 359240 49774
rect 359188 49710 359240 49716
rect 360108 49768 360160 49774
rect 360108 49710 360160 49716
rect 360200 49768 360252 49774
rect 360200 49710 360252 49716
rect 358648 6886 358768 6914
rect 357348 4004 357400 4010
rect 357348 3946 357400 3952
rect 358648 3806 358676 6886
rect 358728 4072 358780 4078
rect 358728 4014 358780 4020
rect 358636 3800 358688 3806
rect 358636 3742 358688 3748
rect 357532 3732 357584 3738
rect 357532 3674 357584 3680
rect 357256 3664 357308 3670
rect 357256 3606 357308 3612
rect 355968 3528 356020 3534
rect 355968 3470 356020 3476
rect 356336 2984 356388 2990
rect 356336 2926 356388 2932
rect 356348 480 356376 2926
rect 357544 480 357572 3674
rect 358740 480 358768 4014
rect 360120 3874 360148 49710
rect 361120 3936 361172 3942
rect 361120 3878 361172 3884
rect 359924 3868 359976 3874
rect 359924 3810 359976 3816
rect 360108 3868 360160 3874
rect 360108 3810 360160 3816
rect 359936 480 359964 3810
rect 361132 480 361160 3878
rect 361408 3466 361436 53094
rect 361488 49768 361540 49774
rect 361488 49710 361540 49716
rect 361500 3738 361528 49710
rect 362880 3942 362908 53094
rect 363248 49774 363276 53108
rect 363236 49768 363288 49774
rect 363236 49710 363288 49716
rect 364156 49768 364208 49774
rect 364156 49710 364208 49716
rect 362868 3936 362920 3942
rect 362868 3878 362920 3884
rect 361488 3732 361540 3738
rect 361488 3674 361540 3680
rect 364168 3602 364196 49710
rect 362316 3596 362368 3602
rect 362316 3538 362368 3544
rect 364156 3596 364208 3602
rect 364156 3538 364208 3544
rect 361396 3460 361448 3466
rect 361396 3402 361448 3408
rect 362328 480 362356 3538
rect 364260 3534 364288 53108
rect 365286 53094 365668 53122
rect 366298 53094 367048 53122
rect 365640 4146 365668 53094
rect 365628 4140 365680 4146
rect 365628 4082 365680 4088
rect 367020 4078 367048 53094
rect 367296 49774 367324 53108
rect 368322 53094 368428 53122
rect 369334 53094 369808 53122
rect 367284 49768 367336 49774
rect 367284 49710 367336 49716
rect 368296 49768 368348 49774
rect 368296 49710 368348 49716
rect 367008 4072 367060 4078
rect 367008 4014 367060 4020
rect 364616 4004 364668 4010
rect 364616 3946 364668 3952
rect 363512 3528 363564 3534
rect 363512 3470 363564 3476
rect 364248 3528 364300 3534
rect 364248 3470 364300 3476
rect 363524 480 363552 3470
rect 364628 480 364656 3946
rect 368204 3868 368256 3874
rect 368204 3810 368256 3816
rect 367008 3800 367060 3806
rect 367008 3742 367060 3748
rect 365812 3664 365864 3670
rect 365812 3606 365864 3612
rect 365824 480 365852 3606
rect 367020 480 367048 3742
rect 368216 480 368244 3810
rect 368308 3806 368336 49710
rect 368296 3800 368348 3806
rect 368296 3742 368348 3748
rect 368400 3670 368428 53094
rect 369780 3738 369808 53094
rect 370332 49774 370360 53108
rect 371344 49774 371372 53108
rect 372370 53094 372476 53122
rect 373382 53094 373948 53122
rect 370320 49768 370372 49774
rect 370320 49710 370372 49716
rect 371148 49768 371200 49774
rect 371148 49710 371200 49716
rect 371332 49768 371384 49774
rect 371332 49710 371384 49716
rect 371160 3874 371188 49710
rect 371700 3936 371752 3942
rect 371700 3878 371752 3884
rect 371148 3868 371200 3874
rect 371148 3810 371200 3816
rect 369400 3732 369452 3738
rect 369400 3674 369452 3680
rect 369768 3732 369820 3738
rect 369768 3674 369820 3680
rect 368388 3664 368440 3670
rect 368388 3606 368440 3612
rect 369412 480 369440 3674
rect 370596 3460 370648 3466
rect 370596 3402 370648 3408
rect 370608 480 370636 3402
rect 371712 480 371740 3878
rect 372448 3466 372476 53094
rect 372528 49768 372580 49774
rect 372528 49710 372580 49716
rect 372540 4010 372568 49710
rect 372528 4004 372580 4010
rect 372528 3946 372580 3952
rect 373920 3942 373948 53094
rect 374380 49774 374408 53108
rect 375392 49774 375420 53108
rect 376418 53094 376708 53122
rect 377522 53094 378088 53122
rect 374368 49768 374420 49774
rect 374368 49710 374420 49716
rect 375288 49768 375340 49774
rect 375288 49710 375340 49716
rect 375380 49768 375432 49774
rect 375380 49710 375432 49716
rect 376576 49768 376628 49774
rect 376576 49710 376628 49716
rect 375300 6914 375328 49710
rect 375208 6886 375328 6914
rect 373908 3936 373960 3942
rect 373908 3878 373960 3884
rect 372896 3596 372948 3602
rect 372896 3538 372948 3544
rect 372436 3460 372488 3466
rect 372436 3402 372488 3408
rect 372908 480 372936 3538
rect 374092 3528 374144 3534
rect 374092 3470 374144 3476
rect 374104 480 374132 3470
rect 375208 3398 375236 6886
rect 375288 4140 375340 4146
rect 375288 4082 375340 4088
rect 375196 3392 375248 3398
rect 375196 3334 375248 3340
rect 375300 480 375328 4082
rect 376484 4072 376536 4078
rect 376484 4014 376536 4020
rect 376496 480 376524 4014
rect 376588 3602 376616 49710
rect 376576 3596 376628 3602
rect 376576 3538 376628 3544
rect 376680 3534 376708 53094
rect 378060 4146 378088 53094
rect 378520 49774 378548 53108
rect 379532 49774 379560 53108
rect 380558 53094 380848 53122
rect 381570 53094 382228 53122
rect 378508 49768 378560 49774
rect 378508 49710 378560 49716
rect 379428 49768 379480 49774
rect 379428 49710 379480 49716
rect 379520 49768 379572 49774
rect 379520 49710 379572 49716
rect 380716 49768 380768 49774
rect 380716 49710 380768 49716
rect 378048 4140 378100 4146
rect 378048 4082 378100 4088
rect 377680 3800 377732 3806
rect 377680 3742 377732 3748
rect 376668 3528 376720 3534
rect 376668 3470 376720 3476
rect 377692 480 377720 3742
rect 379440 3670 379468 49710
rect 379980 3732 380032 3738
rect 379980 3674 380032 3680
rect 378876 3664 378928 3670
rect 378876 3606 378928 3612
rect 379428 3664 379480 3670
rect 379428 3606 379480 3612
rect 378888 480 378916 3606
rect 379992 480 380020 3674
rect 380728 3330 380756 49710
rect 380820 3806 380848 53094
rect 382200 4078 382228 53094
rect 382568 49774 382596 53108
rect 382556 49768 382608 49774
rect 382556 49710 382608 49716
rect 383476 49768 383528 49774
rect 383476 49710 383528 49716
rect 382188 4072 382240 4078
rect 382188 4014 382240 4020
rect 383488 4010 383516 49710
rect 382372 4004 382424 4010
rect 382372 3946 382424 3952
rect 383476 4004 383528 4010
rect 383476 3946 383528 3952
rect 381176 3868 381228 3874
rect 381176 3810 381228 3816
rect 380808 3800 380860 3806
rect 380808 3742 380860 3748
rect 380716 3324 380768 3330
rect 380716 3266 380768 3272
rect 381188 480 381216 3810
rect 382384 480 382412 3946
rect 383580 3584 383608 53108
rect 384606 53094 384988 53122
rect 385618 53094 386368 53122
rect 384960 3942 384988 53094
rect 384764 3936 384816 3942
rect 384764 3878 384816 3884
rect 384948 3936 385000 3942
rect 384948 3878 385000 3884
rect 383580 3556 383700 3584
rect 383672 3466 383700 3556
rect 383568 3460 383620 3466
rect 383568 3402 383620 3408
rect 383660 3460 383712 3466
rect 383660 3402 383712 3408
rect 383580 480 383608 3402
rect 384776 480 384804 3878
rect 386340 3874 386368 53094
rect 386616 49774 386644 53108
rect 386604 49768 386656 49774
rect 386604 49710 386656 49716
rect 386328 3868 386380 3874
rect 386328 3810 386380 3816
rect 387628 3602 387656 53108
rect 388654 53094 389128 53122
rect 387708 49768 387760 49774
rect 387708 49710 387760 49716
rect 387156 3596 387208 3602
rect 387156 3538 387208 3544
rect 387616 3596 387668 3602
rect 387616 3538 387668 3544
rect 385960 3392 386012 3398
rect 385960 3334 386012 3340
rect 385972 480 386000 3334
rect 387168 480 387196 3538
rect 387720 3398 387748 49710
rect 389100 3738 389128 53094
rect 389652 49774 389680 53108
rect 390664 49774 390692 53108
rect 391690 53094 391888 53122
rect 392702 53094 393268 53122
rect 389640 49768 389692 49774
rect 389640 49710 389692 49716
rect 390468 49768 390520 49774
rect 390468 49710 390520 49716
rect 390652 49768 390704 49774
rect 390652 49710 390704 49716
rect 391756 49768 391808 49774
rect 391756 49710 391808 49716
rect 389456 4140 389508 4146
rect 389456 4082 389508 4088
rect 389088 3732 389140 3738
rect 389088 3674 389140 3680
rect 388260 3528 388312 3534
rect 388260 3470 388312 3476
rect 387708 3392 387760 3398
rect 387708 3334 387760 3340
rect 388272 480 388300 3470
rect 389468 480 389496 4082
rect 390480 3194 390508 49710
rect 391768 3670 391796 49710
rect 390652 3664 390704 3670
rect 390652 3606 390704 3612
rect 391756 3664 391808 3670
rect 391756 3606 391808 3612
rect 390468 3188 390520 3194
rect 390468 3130 390520 3136
rect 390664 480 390692 3606
rect 391860 3534 391888 53094
rect 393240 3806 393268 53094
rect 393700 49774 393728 53108
rect 394712 49774 394740 53108
rect 395738 53094 396028 53122
rect 396750 53094 397408 53122
rect 393688 49768 393740 49774
rect 393688 49710 393740 49716
rect 394608 49768 394660 49774
rect 394608 49710 394660 49716
rect 394700 49768 394752 49774
rect 394700 49710 394752 49716
rect 395896 49768 395948 49774
rect 395896 49710 395948 49716
rect 394240 4072 394292 4078
rect 394240 4014 394292 4020
rect 393044 3800 393096 3806
rect 393044 3742 393096 3748
rect 393228 3800 393280 3806
rect 393228 3742 393280 3748
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 391848 3324 391900 3330
rect 391848 3266 391900 3272
rect 391860 480 391888 3266
rect 393056 480 393084 3742
rect 394252 480 394280 4014
rect 394620 3126 394648 49710
rect 395344 4004 395396 4010
rect 395344 3946 395396 3952
rect 394608 3120 394660 3126
rect 394608 3062 394660 3068
rect 395356 480 395384 3946
rect 395908 3330 395936 49710
rect 396000 4078 396028 53094
rect 397380 4146 397408 53094
rect 397748 49774 397776 53108
rect 397736 49768 397788 49774
rect 397736 49710 397788 49716
rect 398656 49768 398708 49774
rect 398656 49710 398708 49716
rect 397368 4140 397420 4146
rect 397368 4082 397420 4088
rect 395988 4072 396040 4078
rect 395988 4014 396040 4020
rect 398668 4010 398696 49710
rect 398656 4004 398708 4010
rect 398656 3946 398708 3952
rect 397736 3936 397788 3942
rect 397736 3878 397788 3884
rect 396540 3460 396592 3466
rect 396540 3402 396592 3408
rect 395896 3324 395948 3330
rect 395896 3266 395948 3272
rect 396552 480 396580 3402
rect 397748 480 397776 3878
rect 398760 3466 398788 53108
rect 399786 53094 400168 53122
rect 400140 3942 400168 53094
rect 400784 49774 400812 53108
rect 401888 49774 401916 53108
rect 402808 53094 402914 53122
rect 403926 53094 404308 53122
rect 404938 53094 405688 53122
rect 400772 49768 400824 49774
rect 400772 49710 400824 49716
rect 401508 49768 401560 49774
rect 401508 49710 401560 49716
rect 401876 49768 401928 49774
rect 401876 49710 401928 49716
rect 400128 3936 400180 3942
rect 400128 3878 400180 3884
rect 398932 3868 398984 3874
rect 398932 3810 398984 3816
rect 398748 3460 398800 3466
rect 398748 3402 398800 3408
rect 398944 480 398972 3810
rect 401324 3596 401376 3602
rect 401324 3538 401376 3544
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 401336 480 401364 3538
rect 401520 3398 401548 49710
rect 402520 3732 402572 3738
rect 402520 3674 402572 3680
rect 401508 3392 401560 3398
rect 401508 3334 401560 3340
rect 402532 480 402560 3674
rect 402808 3602 402836 53094
rect 402888 49768 402940 49774
rect 402888 49710 402940 49716
rect 402796 3596 402848 3602
rect 402796 3538 402848 3544
rect 402900 3262 402928 49710
rect 404280 3738 404308 53094
rect 405660 3874 405688 53094
rect 405936 49774 405964 53108
rect 406962 53094 407068 53122
rect 407974 53094 408448 53122
rect 405924 49768 405976 49774
rect 405924 49710 405976 49716
rect 406936 49768 406988 49774
rect 406936 49710 406988 49716
rect 405648 3868 405700 3874
rect 405648 3810 405700 3816
rect 404268 3732 404320 3738
rect 404268 3674 404320 3680
rect 406948 3670 406976 49710
rect 404820 3664 404872 3670
rect 404820 3606 404872 3612
rect 406936 3664 406988 3670
rect 406936 3606 406988 3612
rect 402888 3256 402940 3262
rect 402888 3198 402940 3204
rect 403624 3188 403676 3194
rect 403624 3130 403676 3136
rect 403636 480 403664 3130
rect 404832 480 404860 3606
rect 407040 3534 407068 53094
rect 408420 6914 408448 53094
rect 408972 49774 409000 53108
rect 409984 49774 410012 53108
rect 411010 53094 411208 53122
rect 412022 53094 412588 53122
rect 408960 49768 409012 49774
rect 408960 49710 409012 49716
rect 409788 49768 409840 49774
rect 409788 49710 409840 49716
rect 409972 49768 410024 49774
rect 409972 49710 410024 49716
rect 411076 49768 411128 49774
rect 411076 49710 411128 49716
rect 408328 6886 408448 6914
rect 407212 3800 407264 3806
rect 407212 3742 407264 3748
rect 406016 3528 406068 3534
rect 406016 3470 406068 3476
rect 407028 3528 407080 3534
rect 407028 3470 407080 3476
rect 406028 480 406056 3470
rect 407224 480 407252 3742
rect 408328 3194 408356 6886
rect 409604 3324 409656 3330
rect 409604 3266 409656 3272
rect 408316 3188 408368 3194
rect 408316 3130 408368 3136
rect 408408 3120 408460 3126
rect 408408 3062 408460 3068
rect 408420 480 408448 3062
rect 409616 480 409644 3266
rect 409800 2922 409828 49710
rect 410800 4072 410852 4078
rect 410800 4014 410852 4020
rect 409788 2916 409840 2922
rect 409788 2858 409840 2864
rect 410812 480 410840 4014
rect 411088 3806 411116 49710
rect 411180 4078 411208 53094
rect 411904 4140 411956 4146
rect 411904 4082 411956 4088
rect 411168 4072 411220 4078
rect 411168 4014 411220 4020
rect 411076 3800 411128 3806
rect 411076 3742 411128 3748
rect 411916 480 411944 4082
rect 412560 3330 412588 53094
rect 413020 49774 413048 53108
rect 414032 49774 414060 53108
rect 415058 53094 415256 53122
rect 416070 53094 416728 53122
rect 413008 49768 413060 49774
rect 413008 49710 413060 49716
rect 413928 49768 413980 49774
rect 413928 49710 413980 49716
rect 414020 49768 414072 49774
rect 414020 49710 414072 49716
rect 413100 4004 413152 4010
rect 413100 3946 413152 3952
rect 412548 3324 412600 3330
rect 412548 3266 412600 3272
rect 413112 480 413140 3946
rect 413940 2990 413968 49710
rect 415228 4010 415256 53094
rect 415308 49768 415360 49774
rect 415308 49710 415360 49716
rect 415320 4146 415348 49710
rect 416700 6914 416728 53094
rect 417068 49774 417096 53108
rect 417988 53094 418094 53122
rect 419106 53094 419488 53122
rect 417056 49768 417108 49774
rect 417056 49710 417108 49716
rect 416608 6886 416728 6914
rect 415308 4140 415360 4146
rect 415308 4082 415360 4088
rect 415216 4004 415268 4010
rect 415216 3946 415268 3952
rect 415492 3936 415544 3942
rect 415492 3878 415544 3884
rect 414296 3460 414348 3466
rect 414296 3402 414348 3408
rect 413928 2984 413980 2990
rect 413928 2926 413980 2932
rect 414308 480 414336 3402
rect 415504 480 415532 3878
rect 416608 3058 416636 6886
rect 417988 3466 418016 53094
rect 418068 49768 418120 49774
rect 418068 49710 418120 49716
rect 417976 3460 418028 3466
rect 417976 3402 418028 3408
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416596 3052 416648 3058
rect 416596 2994 416648 3000
rect 416700 480 416728 3334
rect 418080 3262 418108 49710
rect 419460 3942 419488 53094
rect 420104 49774 420132 53108
rect 421116 49774 421144 53108
rect 420092 49768 420144 49774
rect 420092 49710 420144 49716
rect 420828 49768 420880 49774
rect 420828 49710 420880 49716
rect 421104 49768 421156 49774
rect 421104 49710 421156 49716
rect 419448 3936 419500 3942
rect 419448 3878 419500 3884
rect 420184 3732 420236 3738
rect 420184 3674 420236 3680
rect 418988 3596 419040 3602
rect 418988 3538 419040 3544
rect 417884 3256 417936 3262
rect 417884 3198 417936 3204
rect 418068 3256 418120 3262
rect 418068 3198 418120 3204
rect 417896 480 417924 3198
rect 419000 480 419028 3538
rect 420196 480 420224 3674
rect 420840 3194 420868 49710
rect 421380 3868 421432 3874
rect 421380 3810 421432 3816
rect 420828 3188 420880 3194
rect 420828 3130 420880 3136
rect 421392 480 421420 3810
rect 422128 3602 422156 53108
rect 423154 53094 423628 53122
rect 422208 49768 422260 49774
rect 422208 49710 422260 49716
rect 422220 3738 422248 49710
rect 422208 3732 422260 3738
rect 422208 3674 422260 3680
rect 422576 3664 422628 3670
rect 422576 3606 422628 3612
rect 422116 3596 422168 3602
rect 422116 3538 422168 3544
rect 422588 480 422616 3606
rect 423600 3398 423628 53094
rect 424152 49774 424180 53108
rect 425256 49774 425284 53108
rect 426282 53094 426388 53122
rect 427294 53094 427768 53122
rect 424140 49768 424192 49774
rect 424140 49710 424192 49716
rect 424968 49768 425020 49774
rect 424968 49710 425020 49716
rect 425244 49768 425296 49774
rect 425244 49710 425296 49716
rect 426256 49768 426308 49774
rect 426256 49710 426308 49716
rect 424980 3874 425008 49710
rect 424968 3868 425020 3874
rect 424968 3810 425020 3816
rect 426268 3670 426296 49710
rect 426256 3664 426308 3670
rect 426256 3606 426308 3612
rect 426360 3534 426388 53094
rect 427740 3806 427768 53094
rect 428292 49774 428320 53108
rect 429304 49774 429332 53108
rect 430330 53094 430436 53122
rect 431342 53094 431908 53122
rect 428280 49768 428332 49774
rect 428280 49710 428332 49716
rect 429108 49768 429160 49774
rect 429108 49710 429160 49716
rect 429292 49768 429344 49774
rect 429292 49710 429344 49716
rect 429120 4962 429148 49710
rect 429108 4956 429160 4962
rect 429108 4898 429160 4904
rect 430408 4078 430436 53094
rect 430488 49768 430540 49774
rect 430488 49710 430540 49716
rect 428464 4072 428516 4078
rect 428464 4014 428516 4020
rect 430396 4072 430448 4078
rect 430396 4014 430448 4020
rect 427268 3800 427320 3806
rect 427268 3742 427320 3748
rect 427728 3800 427780 3806
rect 427728 3742 427780 3748
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 426348 3528 426400 3534
rect 426348 3470 426400 3476
rect 423588 3392 423640 3398
rect 423588 3334 423640 3340
rect 423784 480 423812 3470
rect 424968 3120 425020 3126
rect 424968 3062 425020 3068
rect 424980 480 425008 3062
rect 426164 2916 426216 2922
rect 426164 2858 426216 2864
rect 426176 480 426204 2858
rect 427280 480 427308 3742
rect 428476 480 428504 4014
rect 429660 3324 429712 3330
rect 429660 3266 429712 3272
rect 429672 480 429700 3266
rect 430500 3126 430528 49710
rect 431880 5030 431908 53094
rect 432340 49774 432368 53108
rect 433352 49774 433380 53108
rect 434364 49842 434392 53108
rect 435390 53094 436048 53122
rect 434352 49836 434404 49842
rect 434352 49778 434404 49784
rect 435364 49836 435416 49842
rect 435364 49778 435416 49784
rect 432328 49768 432380 49774
rect 432328 49710 432380 49716
rect 433248 49768 433300 49774
rect 433248 49710 433300 49716
rect 433340 49768 433392 49774
rect 433340 49710 433392 49716
rect 434628 49768 434680 49774
rect 434628 49710 434680 49716
rect 431868 5024 431920 5030
rect 431868 4966 431920 4972
rect 433260 4146 433288 49710
rect 432052 4140 432104 4146
rect 432052 4082 432104 4088
rect 433248 4140 433300 4146
rect 433248 4082 433300 4088
rect 430488 3120 430540 3126
rect 430488 3062 430540 3068
rect 430856 2984 430908 2990
rect 430856 2926 430908 2932
rect 430868 480 430896 2926
rect 432064 480 432092 4082
rect 433248 4004 433300 4010
rect 433248 3946 433300 3952
rect 433260 480 433288 3946
rect 434640 3330 434668 49710
rect 435376 4826 435404 49778
rect 435364 4820 435416 4826
rect 435364 4762 435416 4768
rect 436020 4010 436048 53094
rect 436388 49774 436416 53108
rect 437308 53094 437414 53122
rect 438426 53094 438808 53122
rect 436376 49768 436428 49774
rect 436376 49710 436428 49716
rect 437308 4894 437336 53094
rect 437388 49768 437440 49774
rect 437388 49710 437440 49716
rect 437296 4888 437348 4894
rect 437296 4830 437348 4836
rect 436008 4004 436060 4010
rect 436008 3946 436060 3952
rect 436744 3460 436796 3466
rect 436744 3402 436796 3408
rect 434628 3324 434680 3330
rect 434628 3266 434680 3272
rect 435548 3256 435600 3262
rect 435548 3198 435600 3204
rect 434444 3052 434496 3058
rect 434444 2994 434496 3000
rect 434456 480 434484 2994
rect 435560 480 435588 3198
rect 436756 480 436784 3402
rect 437400 3262 437428 49710
rect 438780 3942 438808 53094
rect 439424 49774 439452 53108
rect 440436 50386 440464 53108
rect 441462 53094 441568 53122
rect 442474 53094 442948 53122
rect 440424 50380 440476 50386
rect 440424 50322 440476 50328
rect 439412 49768 439464 49774
rect 439412 49710 439464 49716
rect 440148 49768 440200 49774
rect 440148 49710 440200 49716
rect 437940 3936 437992 3942
rect 437940 3878 437992 3884
rect 438768 3936 438820 3942
rect 438768 3878 438820 3884
rect 437388 3256 437440 3262
rect 437388 3198 437440 3204
rect 437952 480 437980 3878
rect 439136 3188 439188 3194
rect 439136 3130 439188 3136
rect 439148 480 439176 3130
rect 440160 2990 440188 49710
rect 441540 3754 441568 53094
rect 440332 3732 440384 3738
rect 441540 3726 441660 3754
rect 442920 3738 442948 53094
rect 443472 49774 443500 53108
rect 444484 49774 444512 53108
rect 445510 53094 445616 53122
rect 446522 53094 447088 53122
rect 443460 49768 443512 49774
rect 443460 49710 443512 49716
rect 444288 49768 444340 49774
rect 444288 49710 444340 49716
rect 444472 49768 444524 49774
rect 444472 49710 444524 49716
rect 443828 3868 443880 3874
rect 443828 3810 443880 3816
rect 440332 3674 440384 3680
rect 440148 2984 440200 2990
rect 440148 2926 440200 2932
rect 440344 480 440372 3674
rect 441632 3602 441660 3726
rect 442908 3732 442960 3738
rect 442908 3674 442960 3680
rect 441528 3596 441580 3602
rect 441528 3538 441580 3544
rect 441620 3596 441672 3602
rect 441620 3538 441672 3544
rect 441540 480 441568 3538
rect 442632 3392 442684 3398
rect 442632 3334 442684 3340
rect 442644 480 442672 3334
rect 443840 480 443868 3810
rect 444300 2922 444328 49710
rect 445024 3664 445076 3670
rect 445024 3606 445076 3612
rect 444288 2916 444340 2922
rect 444288 2858 444340 2864
rect 445036 480 445064 3606
rect 445588 3466 445616 53094
rect 446404 50380 446456 50386
rect 446404 50322 446456 50328
rect 445668 49768 445720 49774
rect 445668 49710 445720 49716
rect 445576 3460 445628 3466
rect 445576 3402 445628 3408
rect 445680 3058 445708 49710
rect 446416 5166 446444 50322
rect 446404 5160 446456 5166
rect 446404 5102 446456 5108
rect 447060 3670 447088 53094
rect 447520 49774 447548 53108
rect 448532 49774 448560 53108
rect 449650 53094 449756 53122
rect 450662 53094 451228 53122
rect 447508 49768 447560 49774
rect 447508 49710 447560 49716
rect 448428 49768 448480 49774
rect 448428 49710 448480 49716
rect 448520 49768 448572 49774
rect 448520 49710 448572 49716
rect 448440 3874 448468 49710
rect 448612 4956 448664 4962
rect 448612 4898 448664 4904
rect 448428 3868 448480 3874
rect 448428 3810 448480 3816
rect 447416 3800 447468 3806
rect 447416 3742 447468 3748
rect 447048 3664 447100 3670
rect 447048 3606 447100 3612
rect 446220 3528 446272 3534
rect 446220 3470 446272 3476
rect 445668 3052 445720 3058
rect 445668 2994 445720 3000
rect 446232 480 446260 3470
rect 447428 480 447456 3742
rect 448624 480 448652 4898
rect 449728 3534 449756 53094
rect 449808 49768 449860 49774
rect 449808 49710 449860 49716
rect 449820 3806 449848 49710
rect 450912 4072 450964 4078
rect 450912 4014 450964 4020
rect 449808 3800 449860 3806
rect 449808 3742 449860 3748
rect 449716 3528 449768 3534
rect 449716 3470 449768 3476
rect 449808 3120 449860 3126
rect 449808 3062 449860 3068
rect 449820 480 449848 3062
rect 450924 480 450952 4014
rect 451200 3126 451228 53094
rect 451660 49842 451688 53108
rect 451648 49836 451700 49842
rect 451648 49778 451700 49784
rect 452672 49774 452700 53108
rect 453698 53094 453988 53122
rect 454710 53094 455368 53122
rect 452660 49768 452712 49774
rect 452660 49710 452712 49716
rect 453856 49768 453908 49774
rect 453856 49710 453908 49716
rect 452108 5024 452160 5030
rect 452108 4966 452160 4972
rect 451188 3120 451240 3126
rect 451188 3062 451240 3068
rect 452120 480 452148 4966
rect 453304 4140 453356 4146
rect 453304 4082 453356 4088
rect 453316 480 453344 4082
rect 453868 3194 453896 49710
rect 453960 3942 453988 53094
rect 454684 49836 454736 49842
rect 454684 49778 454736 49784
rect 453948 3936 454000 3942
rect 453948 3878 454000 3884
rect 454500 3324 454552 3330
rect 454500 3266 454552 3272
rect 453856 3188 453908 3194
rect 453856 3130 453908 3136
rect 454512 480 454540 3266
rect 454696 2854 454724 49778
rect 455340 3398 455368 53094
rect 455708 49774 455736 53108
rect 455696 49768 455748 49774
rect 455696 49710 455748 49716
rect 455696 4820 455748 4826
rect 455696 4762 455748 4768
rect 455328 3392 455380 3398
rect 455328 3334 455380 3340
rect 454684 2848 454736 2854
rect 454684 2790 454736 2796
rect 455708 480 455736 4762
rect 456720 4078 456748 53108
rect 457746 53094 458128 53122
rect 457444 49768 457496 49774
rect 457444 49710 457496 49716
rect 457456 4826 457484 49710
rect 458100 6914 458128 53094
rect 458744 50794 458772 53108
rect 458732 50788 458784 50794
rect 458732 50730 458784 50736
rect 459756 49774 459784 53108
rect 460782 53094 460888 53122
rect 461794 53094 462268 53122
rect 459744 49768 459796 49774
rect 459744 49710 459796 49716
rect 460756 49768 460808 49774
rect 460756 49710 460808 49716
rect 458008 6886 458128 6914
rect 457444 4820 457496 4826
rect 457444 4762 457496 4768
rect 456708 4072 456760 4078
rect 456708 4014 456760 4020
rect 456892 4004 456944 4010
rect 456892 3946 456944 3952
rect 456904 480 456932 3946
rect 458008 3330 458036 6886
rect 459192 4888 459244 4894
rect 459192 4830 459244 4836
rect 457996 3324 458048 3330
rect 457996 3266 458048 3272
rect 458088 3256 458140 3262
rect 458088 3198 458140 3204
rect 458100 480 458128 3198
rect 459204 480 459232 4830
rect 460768 4146 460796 49710
rect 460388 4140 460440 4146
rect 460388 4082 460440 4088
rect 460756 4140 460808 4146
rect 460756 4082 460808 4088
rect 460400 480 460428 4082
rect 460860 3942 460888 53094
rect 461584 50788 461636 50794
rect 461584 50730 461636 50736
rect 461596 5234 461624 50730
rect 461584 5228 461636 5234
rect 461584 5170 461636 5176
rect 462240 5098 462268 53094
rect 462792 49774 462820 53108
rect 463804 49774 463832 53108
rect 464830 53094 464936 53122
rect 465842 53094 466408 53122
rect 462780 49768 462832 49774
rect 462780 49710 462832 49716
rect 463608 49768 463660 49774
rect 463608 49710 463660 49716
rect 463792 49768 463844 49774
rect 463792 49710 463844 49716
rect 462780 5160 462832 5166
rect 462780 5102 462832 5108
rect 462228 5092 462280 5098
rect 462228 5034 462280 5040
rect 460848 3936 460900 3942
rect 460848 3878 460900 3884
rect 461584 2984 461636 2990
rect 461584 2926 461636 2932
rect 461596 480 461624 2926
rect 462792 480 462820 5102
rect 463620 4010 463648 49710
rect 464908 5030 464936 53094
rect 464988 49768 465040 49774
rect 464988 49710 465040 49716
rect 464896 5024 464948 5030
rect 464896 4966 464948 4972
rect 463608 4004 463660 4010
rect 463608 3946 463660 3952
rect 465000 3602 465028 49710
rect 465172 3732 465224 3738
rect 465172 3674 465224 3680
rect 463976 3596 464028 3602
rect 463976 3538 464028 3544
rect 464988 3596 465040 3602
rect 464988 3538 465040 3544
rect 463988 480 464016 3538
rect 465184 480 465212 3674
rect 466380 2990 466408 53094
rect 466840 49774 466868 53108
rect 467852 49774 467880 53108
rect 468878 53094 469168 53122
rect 469890 53094 470548 53122
rect 466828 49768 466880 49774
rect 466828 49710 466880 49716
rect 467748 49768 467800 49774
rect 467748 49710 467800 49716
rect 467840 49768 467892 49774
rect 467840 49710 467892 49716
rect 469036 49768 469088 49774
rect 469036 49710 469088 49716
rect 467760 3738 467788 49710
rect 469048 4962 469076 49710
rect 469036 4956 469088 4962
rect 469036 4898 469088 4904
rect 467748 3732 467800 3738
rect 467748 3674 467800 3680
rect 469140 3466 469168 53094
rect 470520 3670 470548 53094
rect 470888 49774 470916 53108
rect 470876 49768 470928 49774
rect 470876 49710 470928 49716
rect 471796 49768 471848 49774
rect 471796 49710 471848 49716
rect 471808 4894 471836 49710
rect 471796 4888 471848 4894
rect 471796 4830 471848 4836
rect 471900 3874 471928 53108
rect 473018 53094 473308 53122
rect 471060 3868 471112 3874
rect 471060 3810 471112 3816
rect 471888 3868 471940 3874
rect 471888 3810 471940 3816
rect 469864 3664 469916 3670
rect 469864 3606 469916 3612
rect 470508 3664 470560 3670
rect 470508 3606 470560 3612
rect 468668 3460 468720 3466
rect 468668 3402 468720 3408
rect 469128 3460 469180 3466
rect 469128 3402 469180 3408
rect 467472 3052 467524 3058
rect 467472 2994 467524 3000
rect 466368 2984 466420 2990
rect 466368 2926 466420 2932
rect 466276 2916 466328 2922
rect 466276 2858 466328 2864
rect 466288 480 466316 2858
rect 467484 480 467512 2994
rect 468680 480 468708 3402
rect 469876 480 469904 3606
rect 471072 480 471100 3810
rect 472256 3800 472308 3806
rect 472256 3742 472308 3748
rect 472268 480 472296 3742
rect 473280 3058 473308 53094
rect 474016 50386 474044 53108
rect 474004 50380 474056 50386
rect 474004 50322 474056 50328
rect 475028 49774 475056 53108
rect 475016 49768 475068 49774
rect 475016 49710 475068 49716
rect 475936 49768 475988 49774
rect 475936 49710 475988 49716
rect 475948 3806 475976 49710
rect 475936 3800 475988 3806
rect 475936 3742 475988 3748
rect 476040 3534 476068 53108
rect 477052 50794 477080 53108
rect 477040 50788 477092 50794
rect 477040 50730 477092 50736
rect 478064 49774 478092 53108
rect 479076 49774 479104 53108
rect 478052 49768 478104 49774
rect 478052 49710 478104 49716
rect 478788 49768 478840 49774
rect 478788 49710 478840 49716
rect 479064 49768 479116 49774
rect 479064 49710 479116 49716
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 476028 3528 476080 3534
rect 476028 3470 476080 3476
rect 473268 3052 473320 3058
rect 473268 2994 473320 3000
rect 473464 480 473492 3470
rect 478800 3398 478828 49710
rect 480088 5166 480116 53108
rect 481114 53094 481588 53122
rect 480168 49768 480220 49774
rect 480168 49710 480220 49716
rect 480076 5160 480128 5166
rect 480076 5102 480128 5108
rect 478144 3392 478196 3398
rect 478144 3334 478196 3340
rect 478788 3392 478840 3398
rect 478788 3334 478840 3340
rect 476948 3188 477000 3194
rect 476948 3130 477000 3136
rect 474556 3120 474608 3126
rect 474556 3062 474608 3068
rect 474568 480 474596 3062
rect 475752 2848 475804 2854
rect 475752 2790 475804 2796
rect 475764 480 475792 2790
rect 476960 480 476988 3130
rect 478156 480 478184 3334
rect 479340 3324 479392 3330
rect 479340 3266 479392 3272
rect 479352 480 479380 3266
rect 480180 3126 480208 49710
rect 480536 4820 480588 4826
rect 480536 4762 480588 4768
rect 480168 3120 480220 3126
rect 480168 3062 480220 3068
rect 480548 480 480576 4762
rect 481560 3330 481588 53094
rect 482112 49774 482140 53108
rect 482284 50788 482336 50794
rect 482284 50730 482336 50736
rect 482100 49768 482152 49774
rect 482100 49710 482152 49716
rect 482296 5302 482324 50730
rect 483124 49774 483152 53108
rect 484150 53094 484348 53122
rect 485162 53094 485728 53122
rect 482928 49768 482980 49774
rect 482928 49710 482980 49716
rect 483112 49768 483164 49774
rect 483112 49710 483164 49716
rect 484216 49768 484268 49774
rect 484216 49710 484268 49716
rect 482284 5296 482336 5302
rect 482284 5238 482336 5244
rect 481732 4072 481784 4078
rect 481732 4014 481784 4020
rect 481548 3324 481600 3330
rect 481548 3266 481600 3272
rect 481744 480 481772 4014
rect 482836 3256 482888 3262
rect 482836 3198 482888 3204
rect 482848 480 482876 3198
rect 482940 3194 482968 49710
rect 484032 5228 484084 5234
rect 484032 5170 484084 5176
rect 482928 3188 482980 3194
rect 482928 3130 482980 3136
rect 484044 480 484072 5170
rect 484228 4826 484256 49710
rect 484216 4820 484268 4826
rect 484216 4762 484268 4768
rect 484320 4078 484348 53094
rect 485700 4146 485728 53094
rect 486160 49774 486188 53108
rect 487172 49774 487200 53108
rect 488184 50454 488212 53108
rect 489210 53094 489868 53122
rect 488172 50448 488224 50454
rect 488172 50390 488224 50396
rect 486148 49768 486200 49774
rect 486148 49710 486200 49716
rect 487068 49768 487120 49774
rect 487068 49710 487120 49716
rect 487160 49768 487212 49774
rect 487160 49710 487212 49716
rect 488448 49768 488500 49774
rect 488448 49710 488500 49716
rect 487080 5234 487108 49710
rect 487068 5228 487120 5234
rect 487068 5170 487120 5176
rect 487620 5092 487672 5098
rect 487620 5034 487672 5040
rect 485228 4140 485280 4146
rect 485228 4082 485280 4088
rect 485688 4140 485740 4146
rect 485688 4082 485740 4088
rect 484308 4072 484360 4078
rect 484308 4014 484360 4020
rect 485240 480 485268 4082
rect 486424 3936 486476 3942
rect 486424 3878 486476 3884
rect 486436 480 486464 3878
rect 487632 480 487660 5034
rect 488460 3262 488488 49710
rect 489840 5098 489868 53094
rect 490208 49774 490236 53108
rect 490196 49768 490248 49774
rect 490196 49710 490248 49716
rect 491116 49768 491168 49774
rect 491116 49710 491168 49716
rect 489828 5092 489880 5098
rect 489828 5034 489880 5040
rect 491024 5024 491076 5030
rect 491024 4966 491076 4972
rect 488816 4004 488868 4010
rect 488816 3946 488868 3952
rect 488448 3256 488500 3262
rect 488448 3198 488500 3204
rect 488828 480 488856 3946
rect 489920 3596 489972 3602
rect 489920 3538 489972 3544
rect 489932 480 489960 3538
rect 491036 2530 491064 4966
rect 491128 3942 491156 49710
rect 491116 3936 491168 3942
rect 491116 3878 491168 3884
rect 491220 3602 491248 53108
rect 492232 50658 492260 53108
rect 493258 53094 494008 53122
rect 492220 50652 492272 50658
rect 492220 50594 492272 50600
rect 493324 50380 493376 50386
rect 493324 50322 493376 50328
rect 493336 4486 493364 50322
rect 493324 4480 493376 4486
rect 493324 4422 493376 4428
rect 493980 4010 494008 53094
rect 494256 50522 494284 53108
rect 495268 50590 495296 53108
rect 496294 53094 496768 53122
rect 495256 50584 495308 50590
rect 495256 50526 495308 50532
rect 494244 50516 494296 50522
rect 494244 50458 494296 50464
rect 494704 4956 494756 4962
rect 494704 4898 494756 4904
rect 493968 4004 494020 4010
rect 493968 3946 494020 3952
rect 493508 3732 493560 3738
rect 493508 3674 493560 3680
rect 491208 3596 491260 3602
rect 491208 3538 491260 3544
rect 492312 2984 492364 2990
rect 492312 2926 492364 2932
rect 491036 2502 491156 2530
rect 491128 480 491156 2502
rect 492324 480 492352 2926
rect 493520 480 493548 3674
rect 494716 480 494744 4898
rect 496740 3738 496768 53094
rect 497384 49774 497412 53108
rect 498396 50454 498424 53108
rect 499422 53094 499528 53122
rect 500434 53094 500908 53122
rect 497464 50448 497516 50454
rect 497464 50390 497516 50396
rect 498384 50448 498436 50454
rect 498384 50390 498436 50396
rect 497372 49768 497424 49774
rect 497372 49710 497424 49716
rect 496728 3732 496780 3738
rect 496728 3674 496780 3680
rect 497096 3664 497148 3670
rect 497096 3606 497148 3612
rect 495900 3460 495952 3466
rect 495900 3402 495952 3408
rect 495912 480 495940 3402
rect 497108 480 497136 3606
rect 497476 2990 497504 50390
rect 498108 49768 498160 49774
rect 498108 49710 498160 49716
rect 498120 3670 498148 49710
rect 498200 4888 498252 4894
rect 498200 4830 498252 4836
rect 498108 3664 498160 3670
rect 498108 3606 498160 3612
rect 497464 2984 497516 2990
rect 497464 2926 497516 2932
rect 498212 480 498240 4830
rect 499396 3868 499448 3874
rect 499396 3810 499448 3816
rect 499408 480 499436 3810
rect 499500 3466 499528 53094
rect 500224 50652 500276 50658
rect 500224 50594 500276 50600
rect 500236 5370 500264 50594
rect 500224 5364 500276 5370
rect 500224 5306 500276 5312
rect 500880 3874 500908 53094
rect 501432 49774 501460 53108
rect 502444 49774 502472 53108
rect 503456 50386 503484 53108
rect 504482 53094 505048 53122
rect 504364 50584 504416 50590
rect 504364 50526 504416 50532
rect 503444 50380 503496 50386
rect 503444 50322 503496 50328
rect 501420 49768 501472 49774
rect 501420 49710 501472 49716
rect 502248 49768 502300 49774
rect 502248 49710 502300 49716
rect 502432 49768 502484 49774
rect 502432 49710 502484 49716
rect 503628 49768 503680 49774
rect 503628 49710 503680 49716
rect 502260 5030 502288 49710
rect 502248 5024 502300 5030
rect 502248 4966 502300 4972
rect 501788 4480 501840 4486
rect 501788 4422 501840 4428
rect 500868 3868 500920 3874
rect 500868 3810 500920 3816
rect 499488 3460 499540 3466
rect 499488 3402 499540 3408
rect 500592 3052 500644 3058
rect 500592 2994 500644 3000
rect 500604 480 500632 2994
rect 501800 480 501828 4422
rect 503640 3806 503668 49710
rect 504376 5438 504404 50526
rect 504364 5432 504416 5438
rect 504364 5374 504416 5380
rect 505020 4962 505048 53094
rect 505480 49774 505508 53108
rect 506492 50862 506520 53108
rect 507518 53094 507808 53122
rect 508530 53094 509188 53122
rect 506480 50856 506532 50862
rect 506480 50798 506532 50804
rect 505468 49768 505520 49774
rect 505468 49710 505520 49716
rect 506388 49768 506440 49774
rect 506388 49710 506440 49716
rect 505376 5296 505428 5302
rect 505376 5238 505428 5244
rect 505008 4956 505060 4962
rect 505008 4898 505060 4904
rect 502984 3800 503036 3806
rect 502984 3742 503036 3748
rect 503628 3800 503680 3806
rect 503628 3742 503680 3748
rect 502996 480 503024 3742
rect 504180 3528 504232 3534
rect 504180 3470 504232 3476
rect 504192 480 504220 3470
rect 505388 480 505416 5238
rect 506400 3534 506428 49710
rect 507780 4894 507808 53094
rect 508872 5160 508924 5166
rect 508872 5102 508924 5108
rect 507768 4888 507820 4894
rect 507768 4830 507820 4836
rect 506388 3528 506440 3534
rect 506388 3470 506440 3476
rect 506480 3392 506532 3398
rect 506480 3334 506532 3340
rect 506492 480 506520 3334
rect 507676 3120 507728 3126
rect 507676 3062 507728 3068
rect 507688 480 507716 3062
rect 508884 480 508912 5102
rect 509160 3058 509188 53094
rect 509528 50930 509556 53108
rect 510540 50998 510568 53108
rect 511566 53094 511948 53122
rect 512578 53094 513328 53122
rect 510528 50992 510580 50998
rect 510528 50934 510580 50940
rect 509516 50924 509568 50930
rect 509516 50866 509568 50872
rect 511920 3398 511948 53094
rect 512460 4820 512512 4826
rect 512460 4762 512512 4768
rect 511908 3392 511960 3398
rect 511908 3334 511960 3340
rect 510068 3324 510120 3330
rect 510068 3266 510120 3272
rect 509148 3052 509200 3058
rect 509148 2994 509200 3000
rect 510080 480 510108 3266
rect 511264 3188 511316 3194
rect 511264 3130 511316 3136
rect 511276 480 511304 3130
rect 512472 480 512500 4762
rect 513300 3126 513328 53094
rect 513576 49910 513604 53108
rect 514602 53094 514708 53122
rect 515614 53094 516088 53122
rect 513564 49904 513616 49910
rect 513564 49846 513616 49852
rect 513564 4072 513616 4078
rect 513564 4014 513616 4020
rect 513288 3120 513340 3126
rect 513288 3062 513340 3068
rect 513576 480 513604 4014
rect 514680 3330 514708 53094
rect 515404 50516 515456 50522
rect 515404 50458 515456 50464
rect 515416 4146 515444 50458
rect 515956 5228 516008 5234
rect 515956 5170 516008 5176
rect 514760 4140 514812 4146
rect 514760 4082 514812 4088
rect 515404 4140 515456 4146
rect 515404 4082 515456 4088
rect 514668 3324 514720 3330
rect 514668 3266 514720 3272
rect 514772 480 514800 4082
rect 515968 480 515996 5170
rect 516060 3194 516088 53094
rect 516612 50794 516640 53108
rect 516600 50788 516652 50794
rect 516600 50730 516652 50736
rect 517624 49774 517652 53108
rect 518650 53094 518848 53122
rect 517612 49768 517664 49774
rect 517612 49710 517664 49716
rect 518716 49768 518768 49774
rect 518716 49710 518768 49716
rect 518728 4826 518756 49710
rect 518716 4820 518768 4826
rect 518716 4762 518768 4768
rect 518820 4078 518848 53094
rect 519648 50590 519676 53108
rect 519636 50584 519688 50590
rect 519636 50526 519688 50532
rect 519544 49904 519596 49910
rect 519544 49846 519596 49852
rect 519556 5098 519584 49846
rect 520752 49774 520780 53108
rect 520924 50788 520976 50794
rect 520924 50730 520976 50736
rect 520740 49768 520792 49774
rect 520740 49710 520792 49716
rect 520936 6186 520964 50730
rect 521764 49774 521792 53108
rect 522776 50794 522804 53108
rect 523802 53094 524368 53122
rect 522764 50788 522816 50794
rect 522764 50730 522816 50736
rect 521568 49768 521620 49774
rect 521568 49710 521620 49716
rect 521752 49768 521804 49774
rect 521752 49710 521804 49716
rect 522948 49768 523000 49774
rect 522948 49710 523000 49716
rect 520924 6180 520976 6186
rect 520924 6122 520976 6128
rect 519452 5092 519504 5098
rect 519452 5034 519504 5040
rect 519544 5092 519596 5098
rect 519544 5034 519596 5040
rect 518808 4072 518860 4078
rect 518808 4014 518860 4020
rect 517152 3256 517204 3262
rect 517152 3198 517204 3204
rect 516048 3188 516100 3194
rect 516048 3130 516100 3136
rect 517164 480 517192 3198
rect 518348 2984 518400 2990
rect 518348 2926 518400 2932
rect 518360 480 518388 2926
rect 519464 2530 519492 5034
rect 521580 3942 521608 49710
rect 520740 3936 520792 3942
rect 520740 3878 520792 3884
rect 521568 3936 521620 3942
rect 521568 3878 521620 3884
rect 519464 2502 519584 2530
rect 519556 480 519584 2502
rect 520752 480 520780 3878
rect 521844 3596 521896 3602
rect 521844 3538 521896 3544
rect 521856 480 521884 3538
rect 522960 3262 522988 49710
rect 523040 5364 523092 5370
rect 523040 5306 523092 5312
rect 522948 3256 523000 3262
rect 522948 3198 523000 3204
rect 523052 480 523080 5306
rect 524340 4010 524368 53094
rect 524800 49774 524828 53108
rect 525812 50726 525840 53108
rect 526838 53094 527128 53122
rect 525800 50720 525852 50726
rect 525800 50662 525852 50668
rect 525064 50448 525116 50454
rect 525064 50390 525116 50396
rect 524788 49768 524840 49774
rect 524788 49710 524840 49716
rect 525076 4690 525104 50390
rect 525708 49768 525760 49774
rect 525708 49710 525760 49716
rect 525064 4684 525116 4690
rect 525064 4626 525116 4632
rect 525720 4146 525748 49710
rect 526628 5432 526680 5438
rect 526628 5374 526680 5380
rect 525432 4140 525484 4146
rect 525432 4082 525484 4088
rect 525708 4140 525760 4146
rect 525708 4082 525760 4088
rect 524236 4004 524288 4010
rect 524236 3946 524288 3952
rect 524328 4004 524380 4010
rect 524328 3946 524380 3952
rect 524248 480 524276 3946
rect 525444 480 525472 4082
rect 526640 480 526668 5374
rect 527100 3602 527128 53094
rect 527836 50318 527864 53108
rect 528848 50658 528876 53108
rect 528836 50652 528888 50658
rect 528836 50594 528888 50600
rect 527824 50312 527876 50318
rect 527824 50254 527876 50260
rect 527824 3732 527876 3738
rect 527824 3674 527876 3680
rect 527088 3596 527140 3602
rect 527088 3538 527140 3544
rect 527836 480 527864 3674
rect 529860 3670 529888 53108
rect 530872 51066 530900 53108
rect 530860 51060 530912 51066
rect 530860 51002 530912 51008
rect 530584 50380 530636 50386
rect 530584 50322 530636 50328
rect 530124 4684 530176 4690
rect 530124 4626 530176 4632
rect 529020 3664 529072 3670
rect 529020 3606 529072 3612
rect 529848 3664 529900 3670
rect 529848 3606 529900 3612
rect 529032 480 529060 3606
rect 530136 480 530164 4626
rect 530596 3466 530624 50322
rect 531884 50250 531912 53108
rect 531872 50244 531924 50250
rect 531872 50186 531924 50192
rect 532896 49774 532924 53108
rect 533908 50182 533936 53108
rect 534920 50386 534948 53108
rect 534908 50380 534960 50386
rect 534908 50322 534960 50328
rect 533896 50176 533948 50182
rect 533896 50118 533948 50124
rect 535932 49774 535960 53108
rect 536104 50992 536156 50998
rect 536104 50934 536156 50940
rect 532884 49768 532936 49774
rect 532884 49710 532936 49716
rect 533988 49768 534040 49774
rect 533988 49710 534040 49716
rect 535920 49768 535972 49774
rect 535920 49710 535972 49716
rect 533712 5024 533764 5030
rect 533712 4966 533764 4972
rect 532516 3868 532568 3874
rect 532516 3810 532568 3816
rect 530584 3460 530636 3466
rect 530584 3402 530636 3408
rect 531320 2984 531372 2990
rect 531320 2926 531372 2932
rect 531332 480 531360 2926
rect 532528 480 532556 3810
rect 533724 480 533752 4966
rect 534000 3738 534028 49710
rect 536116 5030 536144 50934
rect 536944 49774 536972 53108
rect 537956 50454 537984 53108
rect 538982 53094 539548 53122
rect 537944 50448 537996 50454
rect 537944 50390 537996 50396
rect 536748 49768 536800 49774
rect 536748 49710 536800 49716
rect 536932 49768 536984 49774
rect 536932 49710 536984 49716
rect 538128 49768 538180 49774
rect 538128 49710 538180 49716
rect 536104 5024 536156 5030
rect 536104 4966 536156 4972
rect 536760 3806 536788 49710
rect 537208 4956 537260 4962
rect 537208 4898 537260 4904
rect 534908 3800 534960 3806
rect 534908 3742 534960 3748
rect 536748 3800 536800 3806
rect 536748 3742 536800 3748
rect 533988 3732 534040 3738
rect 533988 3674 534040 3680
rect 534920 480 534948 3742
rect 536104 3460 536156 3466
rect 536104 3402 536156 3408
rect 536116 480 536144 3402
rect 537220 480 537248 4898
rect 538140 3874 538168 49710
rect 538128 3868 538180 3874
rect 538128 3810 538180 3816
rect 539520 3534 539548 53094
rect 539600 50516 539652 50522
rect 539600 50458 539652 50464
rect 538404 3528 538456 3534
rect 538404 3470 538456 3476
rect 539508 3528 539560 3534
rect 539508 3470 539560 3476
rect 538416 480 538444 3470
rect 539612 480 539640 50458
rect 539980 49774 540008 53108
rect 540244 50312 540296 50318
rect 540244 50254 540296 50260
rect 539968 49768 540020 49774
rect 539968 49710 540020 49716
rect 540256 2990 540284 50254
rect 540992 49910 541020 53108
rect 542018 53094 542308 53122
rect 540980 49904 541032 49910
rect 540980 49846 541032 49852
rect 540796 4888 540848 4894
rect 540796 4830 540848 4836
rect 540244 2984 540296 2990
rect 540244 2926 540296 2932
rect 540808 480 540836 4830
rect 542280 3058 542308 53094
rect 542360 50924 542412 50930
rect 542360 50866 542412 50872
rect 542372 16574 542400 50866
rect 543016 50862 543044 53108
rect 544384 51060 544436 51066
rect 544384 51002 544436 51008
rect 543004 50856 543056 50862
rect 543004 50798 543056 50804
rect 544396 16574 544424 51002
rect 548524 50856 548576 50862
rect 548524 50798 548576 50804
rect 545764 50176 545816 50182
rect 545764 50118 545816 50124
rect 542372 16546 542768 16574
rect 544396 16546 544516 16574
rect 541992 3052 542044 3058
rect 541992 2994 542044 3000
rect 542268 3052 542320 3058
rect 542268 2994 542320 3000
rect 542004 480 542032 2994
rect 542740 490 542768 16546
rect 544384 5024 544436 5030
rect 544384 4966 544436 4972
rect 543016 598 543228 626
rect 543016 490 543044 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 462 543044 490
rect 543200 480 543228 598
rect 544396 480 544424 4966
rect 544488 2854 544516 16546
rect 545488 3392 545540 3398
rect 545488 3334 545540 3340
rect 544476 2848 544528 2854
rect 544476 2790 544528 2796
rect 545500 480 545528 3334
rect 545776 2922 545804 50118
rect 547144 49768 547196 49774
rect 547144 49710 547196 49716
rect 547156 3126 547184 49710
rect 547880 5092 547932 5098
rect 547880 5034 547932 5040
rect 546684 3120 546736 3126
rect 546684 3062 546736 3068
rect 547144 3120 547196 3126
rect 547144 3062 547196 3068
rect 545764 2916 545816 2922
rect 545764 2858 545816 2864
rect 546696 480 546724 3062
rect 547892 480 547920 5034
rect 548536 3398 548564 50798
rect 548616 49904 548668 49910
rect 548616 49846 548668 49852
rect 548628 4078 548656 49846
rect 551296 6866 551324 655551
rect 551388 431934 551416 657834
rect 555516 656328 555568 656334
rect 555516 656270 555568 656276
rect 555422 655752 555478 655761
rect 555422 655687 555478 655696
rect 554044 655308 554096 655314
rect 554044 655250 554096 655256
rect 554056 525774 554084 655250
rect 554044 525768 554096 525774
rect 554044 525710 554096 525716
rect 551376 431928 551428 431934
rect 551376 431870 551428 431876
rect 554780 50584 554832 50590
rect 554780 50526 554832 50532
rect 554792 16574 554820 50526
rect 555436 46918 555464 655687
rect 555528 365702 555556 656270
rect 556804 655580 556856 655586
rect 556804 655522 556856 655528
rect 555606 654120 555662 654129
rect 555606 654055 555662 654064
rect 555620 592006 555648 654055
rect 555608 592000 555660 592006
rect 555608 591942 555660 591948
rect 555516 365696 555568 365702
rect 555516 365638 555568 365644
rect 556816 86970 556844 655522
rect 556908 471986 556936 657902
rect 560942 657384 560998 657393
rect 560942 657319 560998 657328
rect 558184 656940 558236 656946
rect 558184 656882 558236 656888
rect 556896 471980 556948 471986
rect 556896 471922 556948 471928
rect 558196 126954 558224 656882
rect 558368 655376 558420 655382
rect 558368 655318 558420 655324
rect 558276 654832 558328 654838
rect 558276 654774 558328 654780
rect 558288 313274 558316 654774
rect 558380 632058 558408 655318
rect 558368 632052 558420 632058
rect 558368 631994 558420 632000
rect 558276 313268 558328 313274
rect 558276 313210 558328 313216
rect 558184 126948 558236 126954
rect 558184 126890 558236 126896
rect 560956 100706 560984 657319
rect 562416 657280 562468 657286
rect 562416 657222 562468 657228
rect 562322 657112 562378 657121
rect 562322 657047 562378 657056
rect 561036 655784 561088 655790
rect 561036 655726 561088 655732
rect 561048 167006 561076 655726
rect 561126 653304 561182 653313
rect 561126 653239 561182 653248
rect 561140 644434 561168 653239
rect 561128 644428 561180 644434
rect 561128 644370 561180 644376
rect 561036 167000 561088 167006
rect 561036 166942 561088 166948
rect 560944 100700 560996 100706
rect 560944 100642 560996 100648
rect 556804 86964 556856 86970
rect 556804 86906 556856 86912
rect 562336 60722 562364 657047
rect 562428 206990 562456 657222
rect 565084 655920 565136 655926
rect 565084 655862 565136 655868
rect 565096 245614 565124 655862
rect 565188 578202 565216 658174
rect 565176 578196 565228 578202
rect 565176 578138 565228 578144
rect 565084 245608 565136 245614
rect 565084 245550 565136 245556
rect 562416 206984 562468 206990
rect 562416 206926 562468 206932
rect 562324 60716 562376 60722
rect 562324 60658 562376 60664
rect 556804 50788 556856 50794
rect 556804 50730 556856 50736
rect 555424 46912 555476 46918
rect 555424 46854 555476 46860
rect 554792 16546 555004 16574
rect 551284 6860 551336 6866
rect 551284 6802 551336 6808
rect 551468 6180 551520 6186
rect 551468 6122 551520 6128
rect 548616 4072 548668 4078
rect 548616 4014 548668 4020
rect 549168 4072 549220 4078
rect 549168 4014 549220 4020
rect 548524 3392 548576 3398
rect 548524 3334 548576 3340
rect 549180 3330 549208 4014
rect 549076 3324 549128 3330
rect 549076 3266 549128 3272
rect 549168 3324 549220 3330
rect 549168 3266 549220 3272
rect 549088 480 549116 3266
rect 550272 3188 550324 3194
rect 550272 3130 550324 3136
rect 550284 480 550312 3130
rect 551480 480 551508 6122
rect 552664 4820 552716 4826
rect 552664 4762 552716 4768
rect 552676 480 552704 4762
rect 553768 3936 553820 3942
rect 553768 3878 553820 3884
rect 553780 480 553808 3878
rect 554976 480 555004 16546
rect 556816 5574 556844 50730
rect 560944 50720 560996 50726
rect 560944 50662 560996 50668
rect 560956 5574 560984 50662
rect 564532 50652 564584 50658
rect 564532 50594 564584 50600
rect 564544 16574 564572 50594
rect 566476 20670 566504 658242
rect 576216 657824 576268 657830
rect 576216 657766 576268 657772
rect 573456 657688 573508 657694
rect 573456 657630 573508 657636
rect 566556 657552 566608 657558
rect 566556 657494 566608 657500
rect 566568 299470 566596 657494
rect 569224 654628 569276 654634
rect 569224 654570 569276 654576
rect 569236 325650 569264 654570
rect 570602 654528 570658 654537
rect 570602 654463 570658 654472
rect 569314 653848 569370 653857
rect 569314 653783 569370 653792
rect 569328 353258 569356 653783
rect 569316 353252 569368 353258
rect 569316 353194 569368 353200
rect 569224 325644 569276 325650
rect 569224 325586 569276 325592
rect 566556 299464 566608 299470
rect 566556 299406 566608 299412
rect 570616 139398 570644 654463
rect 573364 654424 573416 654430
rect 573364 654366 573416 654372
rect 571984 654288 572036 654294
rect 571984 654230 572036 654236
rect 571996 179382 572024 654230
rect 573376 273222 573404 654366
rect 573468 405686 573496 657630
rect 574836 657620 574888 657626
rect 574836 657562 574888 657568
rect 574742 653440 574798 653449
rect 574742 653375 574798 653384
rect 573456 405680 573508 405686
rect 573456 405622 573508 405628
rect 573364 273216 573416 273222
rect 573364 273158 573416 273164
rect 571984 179376 572036 179382
rect 571984 179318 572036 179324
rect 570604 139392 570656 139398
rect 570604 139334 570656 139340
rect 568580 50516 568632 50522
rect 568580 50458 568632 50464
rect 566464 20664 566516 20670
rect 566464 20606 566516 20612
rect 568592 16574 568620 50458
rect 572812 50380 572864 50386
rect 572812 50322 572864 50328
rect 564544 16546 565216 16574
rect 568592 16546 568712 16574
rect 556804 5568 556856 5574
rect 556804 5510 556856 5516
rect 558552 5568 558604 5574
rect 558552 5510 558604 5516
rect 560944 5568 560996 5574
rect 560944 5510 560996 5516
rect 562048 5568 562100 5574
rect 562048 5510 562100 5516
rect 557356 3256 557408 3262
rect 557356 3198 557408 3204
rect 556160 3188 556212 3194
rect 556160 3130 556212 3136
rect 556172 480 556200 3130
rect 557368 480 557396 3198
rect 558564 480 558592 5510
rect 560852 4140 560904 4146
rect 560852 4082 560904 4088
rect 559748 4004 559800 4010
rect 559748 3946 559800 3952
rect 559760 480 559788 3946
rect 560864 480 560892 4082
rect 562060 480 562088 5510
rect 563244 3596 563296 3602
rect 563244 3538 563296 3544
rect 563256 480 563284 3538
rect 564440 2984 564492 2990
rect 564440 2926 564492 2932
rect 564452 480 564480 2926
rect 565188 490 565216 16546
rect 566832 3664 566884 3670
rect 566832 3606 566884 3612
rect 565464 598 565676 626
rect 565464 490 565492 598
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 462 565492 490
rect 565648 480 565676 598
rect 566844 480 566872 3606
rect 568028 2916 568080 2922
rect 568028 2858 568080 2864
rect 568040 480 568068 2858
rect 568684 490 568712 16546
rect 572824 6914 572852 50322
rect 574756 33114 574784 653375
rect 574848 379506 574876 657562
rect 576124 654220 576176 654226
rect 576124 654162 576176 654168
rect 574836 379500 574888 379506
rect 574836 379442 574888 379448
rect 576136 193186 576164 654162
rect 576228 485790 576256 657766
rect 580356 656192 580408 656198
rect 580356 656134 580408 656140
rect 580264 655444 580316 655450
rect 580264 655386 580316 655392
rect 578884 654356 578936 654362
rect 578884 654298 578936 654304
rect 576216 485784 576268 485790
rect 576216 485726 576268 485732
rect 578896 219065 578924 654298
rect 580172 644428 580224 644434
rect 580172 644370 580224 644376
rect 580184 644065 580212 644370
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580172 632052 580224 632058
rect 580172 631994 580224 632000
rect 580184 630873 580212 631994
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580172 618248 580224 618254
rect 580172 618190 580224 618196
rect 580184 617545 580212 618190
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580172 592000 580224 592006
rect 580172 591942 580224 591948
rect 580184 591025 580212 591942
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 579620 578196 579672 578202
rect 579620 578138 579672 578144
rect 579632 577697 579660 578138
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 579896 525768 579948 525774
rect 579896 525710 579948 525716
rect 579908 524521 579936 525710
rect 579894 524512 579950 524521
rect 579894 524447 579950 524456
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 579620 471980 579672 471986
rect 579620 471922 579672 471928
rect 579632 471481 579660 471922
rect 579618 471472 579674 471481
rect 579618 471407 579674 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 579620 431928 579672 431934
rect 579620 431870 579672 431876
rect 579632 431633 579660 431870
rect 579618 431624 579674 431633
rect 579618 431559 579674 431568
rect 579620 405680 579672 405686
rect 579620 405622 579672 405628
rect 579632 404977 579660 405622
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 580276 258913 580304 655386
rect 580368 418305 580396 656134
rect 580354 418296 580410 418305
rect 580354 418231 580410 418240
rect 580262 258904 580318 258913
rect 580262 258839 580318 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 578882 219056 578938 219065
rect 578882 218991 578938 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 576124 193180 576176 193186
rect 576124 193122 576176 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 575480 50448 575532 50454
rect 575480 50390 575532 50396
rect 574744 33108 574796 33114
rect 574744 33050 574796 33056
rect 575492 16574 575520 50390
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 575492 16546 575888 16574
rect 572732 6886 572852 6914
rect 570328 3732 570380 3738
rect 570328 3674 570380 3680
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 3674
rect 571524 3052 571576 3058
rect 571524 2994 571576 3000
rect 571536 480 571564 2994
rect 572732 480 572760 6886
rect 575112 3868 575164 3874
rect 575112 3810 575164 3816
rect 573916 3800 573968 3806
rect 573916 3742 573968 3748
rect 573928 480 573956 3742
rect 575124 480 575152 3810
rect 575860 490 575888 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 577412 3528 577464 3534
rect 577412 3470 577464 3476
rect 576136 598 576348 626
rect 576136 490 576164 598
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 462 576164 490
rect 576320 480 576348 598
rect 577424 480 577452 3470
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 581000 3324 581052 3330
rect 581000 3266 581052 3272
rect 578608 3120 578660 3126
rect 578608 3062 578660 3068
rect 578620 480 578648 3062
rect 581012 480 581040 3266
rect 582208 480 582236 3402
rect 583392 3392 583444 3398
rect 583392 3334 583444 3340
rect 583404 480 583432 3334
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 4802 657464 4858 657520
rect 3422 654200 3478 654256
rect 3330 632032 3386 632088
rect 3146 619112 3202 619168
rect 3054 606056 3110 606112
rect 3330 579944 3386 580000
rect 3330 566888 3386 566944
rect 3330 553832 3386 553888
rect 3330 527856 3386 527912
rect 3146 514800 3202 514856
rect 2962 501744 3018 501800
rect 3238 475632 3294 475688
rect 3054 462576 3110 462632
rect 3330 449520 3386 449576
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 2962 410488 3018 410544
rect 3330 397432 3386 397488
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 2962 267144 3018 267200
rect 3146 254088 3202 254144
rect 3238 241032 3294 241088
rect 3330 214956 3332 214976
rect 3332 214956 3384 214976
rect 3384 214956 3386 214976
rect 3330 214920 3386 214956
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 3514 201864 3570 201920
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 17222 654336 17278 654392
rect 18602 653656 18658 653712
rect 2778 58520 2834 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 21362 653520 21418 653576
rect 33782 655968 33838 656024
rect 35162 655832 35218 655888
rect 36726 653248 36782 653304
rect 40682 654608 40738 654664
rect 39394 653928 39450 653984
rect 45190 655560 45246 655616
rect 80058 657328 80114 657384
rect 62486 657192 62542 657248
rect 58438 655696 58494 655752
rect 66810 657056 66866 657112
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 528098 657464 528154 657520
rect 519358 655968 519414 656024
rect 532514 655832 532570 655888
rect 547142 657192 547198 657248
rect 49514 655016 49570 655072
rect 93490 655016 93546 655072
rect 150254 655016 150310 655072
rect 207570 655016 207626 655072
rect 220910 655016 220966 655072
rect 378506 655016 378562 655072
rect 392122 655016 392178 655072
rect 497002 655016 497058 655072
rect 510250 655016 510306 655072
rect 514758 655016 514814 655072
rect 523590 655016 523646 655072
rect 536838 655016 536894 655072
rect 551282 655560 551338 655616
rect 555422 655696 555478 655752
rect 555606 654064 555662 654120
rect 560942 657328 560998 657384
rect 562322 657056 562378 657112
rect 561126 653248 561182 653304
rect 570602 654472 570658 654528
rect 569314 653792 569370 653848
rect 574742 653384 574798 653440
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 579618 577632 579674 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 537784 580226 537840
rect 579894 524456 579950 524512
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579618 471416 579674 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 579618 431568 579674 431624
rect 579618 404912 579674 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 579618 298696 579674 298752
rect 579894 272176 579950 272232
rect 580354 418240 580410 418296
rect 580262 258848 580318 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 578882 219000 578938 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 4797 657522 4863 657525
rect 528093 657522 528159 657525
rect 4797 657520 528159 657522
rect 4797 657464 4802 657520
rect 4858 657464 528098 657520
rect 528154 657464 528159 657520
rect 4797 657462 528159 657464
rect 4797 657459 4863 657462
rect 528093 657459 528159 657462
rect 80053 657386 80119 657389
rect 560937 657386 561003 657389
rect 80053 657384 561003 657386
rect 80053 657328 80058 657384
rect 80114 657328 560942 657384
rect 560998 657328 561003 657384
rect 80053 657326 561003 657328
rect 80053 657323 80119 657326
rect 560937 657323 561003 657326
rect 62481 657250 62547 657253
rect 547137 657250 547203 657253
rect 62481 657248 547203 657250
rect 62481 657192 62486 657248
rect 62542 657192 547142 657248
rect 547198 657192 547203 657248
rect 583520 657236 584960 657476
rect 62481 657190 547203 657192
rect 62481 657187 62547 657190
rect 547137 657187 547203 657190
rect 66805 657114 66871 657117
rect 562317 657114 562383 657117
rect 66805 657112 562383 657114
rect 66805 657056 66810 657112
rect 66866 657056 562322 657112
rect 562378 657056 562383 657112
rect 66805 657054 562383 657056
rect 66805 657051 66871 657054
rect 562317 657051 562383 657054
rect 33777 656026 33843 656029
rect 519353 656026 519419 656029
rect 33777 656024 519419 656026
rect 33777 655968 33782 656024
rect 33838 655968 519358 656024
rect 519414 655968 519419 656024
rect 33777 655966 519419 655968
rect 33777 655963 33843 655966
rect 519353 655963 519419 655966
rect 35157 655890 35223 655893
rect 532509 655890 532575 655893
rect 35157 655888 532575 655890
rect 35157 655832 35162 655888
rect 35218 655832 532514 655888
rect 532570 655832 532575 655888
rect 35157 655830 532575 655832
rect 35157 655827 35223 655830
rect 532509 655827 532575 655830
rect 58433 655754 58499 655757
rect 555417 655754 555483 655757
rect 58433 655752 555483 655754
rect 58433 655696 58438 655752
rect 58494 655696 555422 655752
rect 555478 655696 555483 655752
rect 58433 655694 555483 655696
rect 58433 655691 58499 655694
rect 555417 655691 555483 655694
rect 45185 655618 45251 655621
rect 551277 655618 551343 655621
rect 45185 655616 551343 655618
rect 45185 655560 45190 655616
rect 45246 655560 551282 655616
rect 551338 655560 551343 655616
rect 45185 655558 551343 655560
rect 45185 655555 45251 655558
rect 551277 655555 551343 655558
rect 49509 655076 49575 655077
rect 49509 655072 49556 655076
rect 49620 655074 49626 655076
rect 93485 655074 93551 655077
rect 150249 655076 150315 655077
rect 98678 655074 98684 655076
rect 49509 655016 49514 655072
rect 49509 655012 49556 655016
rect 49620 655014 49666 655074
rect 93485 655072 98684 655074
rect 93485 655016 93490 655072
rect 93546 655016 98684 655072
rect 93485 655014 98684 655016
rect 49620 655012 49626 655014
rect 49509 655011 49575 655012
rect 93485 655011 93551 655014
rect 98678 655012 98684 655014
rect 98748 655012 98754 655076
rect 150198 655074 150204 655076
rect 150158 655014 150204 655074
rect 150268 655072 150315 655076
rect 150310 655016 150315 655072
rect 150198 655012 150204 655014
rect 150268 655012 150315 655016
rect 150249 655011 150315 655012
rect 207565 655076 207631 655077
rect 207565 655072 207612 655076
rect 207676 655074 207682 655076
rect 220905 655074 220971 655077
rect 221958 655074 221964 655076
rect 207565 655016 207570 655072
rect 207565 655012 207612 655016
rect 207676 655014 207722 655074
rect 220905 655072 221964 655074
rect 220905 655016 220910 655072
rect 220966 655016 221964 655072
rect 220905 655014 221964 655016
rect 207676 655012 207682 655014
rect 207565 655011 207631 655012
rect 220905 655011 220971 655014
rect 221958 655012 221964 655014
rect 222028 655012 222034 655076
rect 376886 655012 376892 655076
rect 376956 655074 376962 655076
rect 378501 655074 378567 655077
rect 376956 655072 378567 655074
rect 376956 655016 378506 655072
rect 378562 655016 378567 655072
rect 376956 655014 378567 655016
rect 376956 655012 376962 655014
rect 378501 655011 378567 655014
rect 392117 655076 392183 655077
rect 392117 655072 392164 655076
rect 392228 655074 392234 655076
rect 496997 655074 497063 655077
rect 392117 655016 392122 655072
rect 392117 655012 392164 655016
rect 392228 655014 392274 655074
rect 489870 655072 497063 655074
rect 489870 655016 497002 655072
rect 497058 655016 497063 655072
rect 489870 655014 497063 655016
rect 392228 655012 392234 655014
rect 392117 655011 392183 655012
rect 222326 654740 222332 654804
rect 222396 654802 222402 654804
rect 231710 654802 231716 654804
rect 222396 654742 231716 654802
rect 222396 654740 222402 654742
rect 231710 654740 231716 654742
rect 231780 654740 231786 654804
rect 231894 654740 231900 654804
rect 231964 654802 231970 654804
rect 241278 654802 241284 654804
rect 231964 654742 241284 654802
rect 231964 654740 231970 654742
rect 241278 654740 241284 654742
rect 241348 654740 241354 654804
rect 241646 654740 241652 654804
rect 241716 654802 241722 654804
rect 251030 654802 251036 654804
rect 241716 654742 251036 654802
rect 241716 654740 241722 654742
rect 251030 654740 251036 654742
rect 251100 654740 251106 654804
rect 251214 654740 251220 654804
rect 251284 654802 251290 654804
rect 260598 654802 260604 654804
rect 251284 654742 260604 654802
rect 251284 654740 251290 654742
rect 260598 654740 260604 654742
rect 260668 654740 260674 654804
rect 260966 654740 260972 654804
rect 261036 654802 261042 654804
rect 270350 654802 270356 654804
rect 261036 654742 270356 654802
rect 261036 654740 261042 654742
rect 270350 654740 270356 654742
rect 270420 654740 270426 654804
rect 270534 654740 270540 654804
rect 270604 654802 270610 654804
rect 279918 654802 279924 654804
rect 270604 654742 279924 654802
rect 270604 654740 270610 654742
rect 279918 654740 279924 654742
rect 279988 654740 279994 654804
rect 280286 654740 280292 654804
rect 280356 654802 280362 654804
rect 289670 654802 289676 654804
rect 280356 654742 289676 654802
rect 280356 654740 280362 654742
rect 289670 654740 289676 654742
rect 289740 654740 289746 654804
rect 289854 654740 289860 654804
rect 289924 654802 289930 654804
rect 299238 654802 299244 654804
rect 289924 654742 299244 654802
rect 289924 654740 289930 654742
rect 299238 654740 299244 654742
rect 299308 654740 299314 654804
rect 299606 654740 299612 654804
rect 299676 654802 299682 654804
rect 308990 654802 308996 654804
rect 299676 654742 308996 654802
rect 299676 654740 299682 654742
rect 308990 654740 308996 654742
rect 309060 654740 309066 654804
rect 309174 654740 309180 654804
rect 309244 654802 309250 654804
rect 318558 654802 318564 654804
rect 309244 654742 318564 654802
rect 309244 654740 309250 654742
rect 318558 654740 318564 654742
rect 318628 654740 318634 654804
rect 318926 654740 318932 654804
rect 318996 654802 319002 654804
rect 328310 654802 328316 654804
rect 318996 654742 328316 654802
rect 318996 654740 319002 654742
rect 328310 654740 328316 654742
rect 328380 654740 328386 654804
rect 328494 654740 328500 654804
rect 328564 654802 328570 654804
rect 337878 654802 337884 654804
rect 328564 654742 337884 654802
rect 328564 654740 328570 654742
rect 337878 654740 337884 654742
rect 337948 654740 337954 654804
rect 338246 654740 338252 654804
rect 338316 654802 338322 654804
rect 347630 654802 347636 654804
rect 338316 654742 347636 654802
rect 338316 654740 338322 654742
rect 347630 654740 347636 654742
rect 347700 654740 347706 654804
rect 347814 654740 347820 654804
rect 347884 654802 347890 654804
rect 357198 654802 357204 654804
rect 347884 654742 357204 654802
rect 347884 654740 347890 654742
rect 357198 654740 357204 654742
rect 357268 654740 357274 654804
rect 357566 654740 357572 654804
rect 357636 654802 357642 654804
rect 366950 654802 366956 654804
rect 357636 654742 366956 654802
rect 357636 654740 357642 654742
rect 366950 654740 366956 654742
rect 367020 654740 367026 654804
rect 367134 654740 367140 654804
rect 367204 654802 367210 654804
rect 376518 654802 376524 654804
rect 367204 654742 376524 654802
rect 367204 654740 367210 654742
rect 376518 654740 376524 654742
rect 376588 654740 376594 654804
rect 40677 654666 40743 654669
rect 489870 654666 489930 655014
rect 496997 655011 497063 655014
rect 504398 655012 504404 655076
rect 504468 655074 504474 655076
rect 510245 655074 510311 655077
rect 504468 655072 510311 655074
rect 504468 655016 510250 655072
rect 510306 655016 510311 655072
rect 504468 655014 510311 655016
rect 504468 655012 504474 655014
rect 510245 655011 510311 655014
rect 512126 655012 512132 655076
rect 512196 655074 512202 655076
rect 514753 655074 514819 655077
rect 523585 655076 523651 655077
rect 536833 655076 536899 655077
rect 523534 655074 523540 655076
rect 512196 655072 514819 655074
rect 512196 655016 514758 655072
rect 514814 655016 514819 655072
rect 512196 655014 514819 655016
rect 523494 655014 523540 655074
rect 523604 655072 523651 655076
rect 536782 655074 536788 655076
rect 523646 655016 523651 655072
rect 512196 655012 512202 655014
rect 514753 655011 514819 655014
rect 523534 655012 523540 655014
rect 523604 655012 523651 655016
rect 536742 655014 536788 655074
rect 536852 655072 536899 655076
rect 536894 655016 536899 655072
rect 536782 655012 536788 655014
rect 536852 655012 536899 655016
rect 523585 655011 523651 655012
rect 536833 655011 536899 655012
rect 40677 654664 489930 654666
rect 40677 654608 40682 654664
rect 40738 654608 489930 654664
rect 40677 654606 489930 654608
rect 40677 654603 40743 654606
rect 98678 654468 98684 654532
rect 98748 654530 98754 654532
rect 570597 654530 570663 654533
rect 98748 654528 570663 654530
rect 98748 654472 570602 654528
rect 570658 654472 570663 654528
rect 98748 654470 570663 654472
rect 98748 654468 98754 654470
rect 570597 654467 570663 654470
rect 17217 654394 17283 654397
rect 504398 654394 504404 654396
rect 17217 654392 504404 654394
rect 17217 654336 17222 654392
rect 17278 654336 504404 654392
rect 17217 654334 504404 654336
rect 17217 654331 17283 654334
rect 504398 654332 504404 654334
rect 504468 654332 504474 654396
rect 3417 654258 3483 654261
rect 512126 654258 512132 654260
rect 3417 654256 512132 654258
rect 3417 654200 3422 654256
rect 3478 654200 512132 654256
rect 3417 654198 512132 654200
rect 3417 654195 3483 654198
rect 512126 654196 512132 654198
rect 512196 654196 512202 654260
rect 207606 654060 207612 654124
rect 207676 654122 207682 654124
rect 555601 654122 555667 654125
rect 207676 654120 555667 654122
rect 207676 654064 555606 654120
rect 555662 654064 555667 654120
rect 207676 654062 555667 654064
rect 207676 654060 207682 654062
rect 555601 654059 555667 654062
rect 39389 653986 39455 653989
rect 392158 653986 392164 653988
rect 39389 653984 392164 653986
rect 39389 653928 39394 653984
rect 39450 653928 392164 653984
rect 39389 653926 392164 653928
rect 39389 653923 39455 653926
rect 392158 653924 392164 653926
rect 392228 653924 392234 653988
rect 150198 653788 150204 653852
rect 150268 653850 150274 653852
rect 569309 653850 569375 653853
rect 150268 653848 569375 653850
rect 150268 653792 569314 653848
rect 569370 653792 569375 653848
rect 150268 653790 569375 653792
rect 150268 653788 150274 653790
rect 569309 653787 569375 653790
rect 18597 653714 18663 653717
rect 523534 653714 523540 653716
rect 18597 653712 523540 653714
rect 18597 653656 18602 653712
rect 18658 653656 523540 653712
rect 18597 653654 523540 653656
rect 18597 653651 18663 653654
rect 523534 653652 523540 653654
rect 523604 653652 523610 653716
rect 21357 653578 21423 653581
rect 536782 653578 536788 653580
rect 21357 653576 536788 653578
rect 21357 653520 21362 653576
rect 21418 653520 536788 653576
rect 21357 653518 536788 653520
rect 21357 653515 21423 653518
rect 536782 653516 536788 653518
rect 536852 653516 536858 653580
rect 49550 653380 49556 653444
rect 49620 653442 49626 653444
rect 574737 653442 574803 653445
rect 49620 653440 574803 653442
rect 49620 653384 574742 653440
rect 574798 653384 574803 653440
rect 49620 653382 574803 653384
rect 49620 653380 49626 653382
rect 574737 653379 574803 653382
rect 36721 653306 36787 653309
rect 222326 653306 222332 653308
rect 36721 653304 222332 653306
rect 36721 653248 36726 653304
rect 36782 653248 222332 653304
rect 36721 653246 222332 653248
rect 36721 653243 36787 653246
rect 222326 653244 222332 653246
rect 222396 653244 222402 653308
rect 222510 653244 222516 653308
rect 222580 653306 222586 653308
rect 561121 653306 561187 653309
rect 222580 653304 561187 653306
rect 222580 653248 561126 653304
rect 561182 653248 561187 653304
rect 222580 653246 561187 653248
rect 222580 653244 222586 653246
rect 561121 653243 561187 653246
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3325 632090 3391 632093
rect -960 632088 3391 632090
rect -960 632032 3330 632088
rect 3386 632032 3391 632088
rect -960 632030 3391 632032
rect -960 631940 480 632030
rect 3325 632027 3391 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3049 606114 3115 606117
rect -960 606112 3115 606114
rect -960 606056 3054 606112
rect 3110 606056 3115 606112
rect -960 606054 3115 606056
rect -960 605964 480 606054
rect 3049 606051 3115 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 579889 524514 579955 524517
rect 583520 524514 584960 524604
rect 579889 524512 584960 524514
rect 579889 524456 579894 524512
rect 579950 524456 584960 524512
rect 579889 524454 584960 524456
rect 579889 524451 579955 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3141 514858 3207 514861
rect -960 514856 3207 514858
rect -960 514800 3146 514856
rect 3202 514800 3207 514856
rect -960 514798 3207 514800
rect -960 514708 480 514798
rect 3141 514795 3207 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2957 501802 3023 501805
rect -960 501800 3023 501802
rect -960 501744 2962 501800
rect 3018 501744 3023 501800
rect -960 501742 3023 501744
rect -960 501652 480 501742
rect 2957 501739 3023 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3233 475690 3299 475693
rect -960 475688 3299 475690
rect -960 475632 3238 475688
rect 3294 475632 3299 475688
rect -960 475630 3299 475632
rect -960 475540 480 475630
rect 3233 475627 3299 475630
rect 579613 471474 579679 471477
rect 583520 471474 584960 471564
rect 579613 471472 584960 471474
rect 579613 471416 579618 471472
rect 579674 471416 584960 471472
rect 579613 471414 584960 471416
rect 579613 471411 579679 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3049 462634 3115 462637
rect -960 462632 3115 462634
rect -960 462576 3054 462632
rect 3110 462576 3115 462632
rect -960 462574 3115 462576
rect -960 462484 480 462574
rect 3049 462571 3115 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579613 431626 579679 431629
rect 583520 431626 584960 431716
rect 579613 431624 584960 431626
rect 579613 431568 579618 431624
rect 579674 431568 584960 431624
rect 579613 431566 584960 431568
rect 579613 431563 579679 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580349 418298 580415 418301
rect 583520 418298 584960 418388
rect 580349 418296 584960 418298
rect 580349 418240 580354 418296
rect 580410 418240 584960 418296
rect 580349 418238 584960 418240
rect 580349 418235 580415 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 579613 404970 579679 404973
rect 583520 404970 584960 405060
rect 579613 404968 584960 404970
rect 579613 404912 579618 404968
rect 579674 404912 584960 404968
rect 579613 404910 584960 404912
rect 579613 404907 579679 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 580257 258906 580323 258909
rect 583520 258906 584960 258996
rect 580257 258904 584960 258906
rect 580257 258848 580262 258904
rect 580318 258848 584960 258904
rect 580257 258846 584960 258848
rect 580257 258843 580323 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 578877 219058 578943 219061
rect 583520 219058 584960 219148
rect 578877 219056 584960 219058
rect 578877 219000 578882 219056
rect 578938 219000 584960 219056
rect 578877 218998 584960 219000
rect 578877 218995 578943 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2773 58578 2839 58581
rect -960 58576 2839 58578
rect -960 58520 2778 58576
rect 2834 58520 2839 58576
rect -960 58518 2839 58520
rect -960 58428 480 58518
rect 2773 58515 2839 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 49556 655072 49620 655076
rect 49556 655016 49570 655072
rect 49570 655016 49620 655072
rect 49556 655012 49620 655016
rect 98684 655012 98748 655076
rect 150204 655072 150268 655076
rect 150204 655016 150254 655072
rect 150254 655016 150268 655072
rect 150204 655012 150268 655016
rect 207612 655072 207676 655076
rect 207612 655016 207626 655072
rect 207626 655016 207676 655072
rect 207612 655012 207676 655016
rect 221964 655012 222028 655076
rect 376892 655012 376956 655076
rect 392164 655072 392228 655076
rect 392164 655016 392178 655072
rect 392178 655016 392228 655072
rect 392164 655012 392228 655016
rect 222332 654740 222396 654804
rect 231716 654740 231780 654804
rect 231900 654740 231964 654804
rect 241284 654740 241348 654804
rect 241652 654740 241716 654804
rect 251036 654740 251100 654804
rect 251220 654740 251284 654804
rect 260604 654740 260668 654804
rect 260972 654740 261036 654804
rect 270356 654740 270420 654804
rect 270540 654740 270604 654804
rect 279924 654740 279988 654804
rect 280292 654740 280356 654804
rect 289676 654740 289740 654804
rect 289860 654740 289924 654804
rect 299244 654740 299308 654804
rect 299612 654740 299676 654804
rect 308996 654740 309060 654804
rect 309180 654740 309244 654804
rect 318564 654740 318628 654804
rect 318932 654740 318996 654804
rect 328316 654740 328380 654804
rect 328500 654740 328564 654804
rect 337884 654740 337948 654804
rect 338252 654740 338316 654804
rect 347636 654740 347700 654804
rect 347820 654740 347884 654804
rect 357204 654740 357268 654804
rect 357572 654740 357636 654804
rect 366956 654740 367020 654804
rect 367140 654740 367204 654804
rect 376524 654740 376588 654804
rect 504404 655012 504468 655076
rect 512132 655012 512196 655076
rect 523540 655072 523604 655076
rect 523540 655016 523590 655072
rect 523590 655016 523604 655072
rect 523540 655012 523604 655016
rect 536788 655072 536852 655076
rect 536788 655016 536838 655072
rect 536838 655016 536852 655072
rect 536788 655012 536852 655016
rect 98684 654468 98748 654532
rect 504404 654332 504468 654396
rect 512132 654196 512196 654260
rect 207612 654060 207676 654124
rect 392164 653924 392228 653988
rect 150204 653788 150268 653852
rect 523540 653652 523604 653716
rect 536788 653516 536852 653580
rect 49556 653380 49620 653444
rect 222332 653244 222396 653308
rect 222516 653244 222580 653308
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 657697 42134 690618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 657697 45854 658338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 657697 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 657697 56414 668898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 657697 60134 672618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 657697 63854 676338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 657697 67574 680058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 657697 74414 686898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 657697 78134 690618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 657697 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 657697 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 657697 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 657697 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 657697 99854 676338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 657697 103574 680058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 657697 110414 686898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 657697 114134 690618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 657697 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 657697 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 657697 128414 668898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 657697 132134 672618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 657697 135854 676338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 657697 139574 680058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 657697 146414 686898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 657697 150134 690618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 657697 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 657697 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 657697 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 657697 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 657697 171854 676338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 657697 175574 680058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 657697 182414 686898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 657697 186134 690618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 657697 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 657697 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 657697 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 657697 204134 672618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 657697 207854 676338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 657697 211574 680058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 657697 218414 686898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 657697 222134 690618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 657697 225854 658338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 657697 229574 662058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 657697 236414 668898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 657697 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 657697 243854 676338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 657697 247574 680058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 657697 254414 686898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 657697 258134 690618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 657697 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 657697 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 657697 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 657697 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 657697 279854 676338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 657697 283574 680058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 657697 290414 686898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 657697 294134 690618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 657697 297854 658338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 657697 301574 662058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 657697 308414 668898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 657697 312134 672618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 657697 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 657697 319574 680058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 657697 326414 686898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 657697 330134 690618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 657697 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 657697 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 657697 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 657697 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 657697 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 657697 355574 680058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 657697 362414 686898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 657697 366134 690618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 657697 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 657697 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 657697 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 657697 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 657697 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 657697 391574 680058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 657697 398414 686898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 657697 402134 690618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 657697 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 657697 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 657697 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 657697 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 657697 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 657697 427574 680058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 657697 434414 686898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 657697 438134 690618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 657697 441854 658338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 657697 445574 662058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 657697 452414 668898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 657697 456134 672618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 657697 459854 676338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 657697 463574 680058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 657697 470414 686898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 657697 474134 690618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 657697 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 657697 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 657697 488414 668898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 657697 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 657697 495854 676338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 657697 499574 680058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 657697 506414 686898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 657697 510134 690618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 657697 513854 658338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 657697 517574 662058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 657697 524414 668898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 657697 528134 672618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 657697 531854 676338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 657697 535574 680058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 657697 542414 686898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 657697 546134 690618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 49555 655076 49621 655077
rect 49555 655012 49556 655076
rect 49620 655012 49621 655076
rect 49555 655011 49621 655012
rect 98683 655076 98749 655077
rect 98683 655012 98684 655076
rect 98748 655012 98749 655076
rect 98683 655011 98749 655012
rect 150203 655076 150269 655077
rect 150203 655012 150204 655076
rect 150268 655012 150269 655076
rect 150203 655011 150269 655012
rect 207611 655076 207677 655077
rect 207611 655012 207612 655076
rect 207676 655012 207677 655076
rect 207611 655011 207677 655012
rect 221963 655076 222029 655077
rect 221963 655012 221964 655076
rect 222028 655012 222029 655076
rect 221963 655011 222029 655012
rect 376891 655076 376957 655077
rect 376891 655012 376892 655076
rect 376956 655012 376957 655076
rect 376891 655011 376957 655012
rect 392163 655076 392229 655077
rect 392163 655012 392164 655076
rect 392228 655012 392229 655076
rect 392163 655011 392229 655012
rect 504403 655076 504469 655077
rect 504403 655012 504404 655076
rect 504468 655012 504469 655076
rect 504403 655011 504469 655012
rect 512131 655076 512197 655077
rect 512131 655012 512132 655076
rect 512196 655012 512197 655076
rect 512131 655011 512197 655012
rect 523539 655076 523605 655077
rect 523539 655012 523540 655076
rect 523604 655012 523605 655076
rect 523539 655011 523605 655012
rect 536787 655076 536853 655077
rect 536787 655012 536788 655076
rect 536852 655012 536853 655076
rect 536787 655011 536853 655012
rect 49558 653445 49618 655011
rect 98686 654533 98746 655011
rect 98683 654532 98749 654533
rect 98683 654468 98684 654532
rect 98748 654468 98749 654532
rect 98683 654467 98749 654468
rect 150206 653853 150266 655011
rect 207614 654125 207674 655011
rect 207611 654124 207677 654125
rect 207611 654060 207612 654124
rect 207676 654060 207677 654124
rect 207611 654059 207677 654060
rect 150203 653852 150269 653853
rect 150203 653788 150204 653852
rect 150268 653788 150269 653852
rect 150203 653787 150269 653788
rect 49555 653444 49621 653445
rect 49555 653380 49556 653444
rect 49620 653380 49621 653444
rect 49555 653379 49621 653380
rect 221966 653170 222026 655011
rect 222331 654804 222397 654805
rect 222331 654740 222332 654804
rect 222396 654740 222397 654804
rect 222331 654739 222397 654740
rect 231715 654804 231781 654805
rect 231715 654740 231716 654804
rect 231780 654740 231781 654804
rect 231715 654739 231781 654740
rect 231899 654804 231965 654805
rect 231899 654740 231900 654804
rect 231964 654740 231965 654804
rect 231899 654739 231965 654740
rect 241283 654804 241349 654805
rect 241283 654740 241284 654804
rect 241348 654740 241349 654804
rect 241283 654739 241349 654740
rect 241651 654804 241717 654805
rect 241651 654740 241652 654804
rect 241716 654740 241717 654804
rect 241651 654739 241717 654740
rect 251035 654804 251101 654805
rect 251035 654740 251036 654804
rect 251100 654740 251101 654804
rect 251035 654739 251101 654740
rect 251219 654804 251285 654805
rect 251219 654740 251220 654804
rect 251284 654740 251285 654804
rect 251219 654739 251285 654740
rect 260603 654804 260669 654805
rect 260603 654740 260604 654804
rect 260668 654740 260669 654804
rect 260603 654739 260669 654740
rect 260971 654804 261037 654805
rect 260971 654740 260972 654804
rect 261036 654740 261037 654804
rect 260971 654739 261037 654740
rect 270355 654804 270421 654805
rect 270355 654740 270356 654804
rect 270420 654740 270421 654804
rect 270355 654739 270421 654740
rect 270539 654804 270605 654805
rect 270539 654740 270540 654804
rect 270604 654740 270605 654804
rect 270539 654739 270605 654740
rect 279923 654804 279989 654805
rect 279923 654740 279924 654804
rect 279988 654740 279989 654804
rect 279923 654739 279989 654740
rect 280291 654804 280357 654805
rect 280291 654740 280292 654804
rect 280356 654740 280357 654804
rect 280291 654739 280357 654740
rect 289675 654804 289741 654805
rect 289675 654740 289676 654804
rect 289740 654740 289741 654804
rect 289675 654739 289741 654740
rect 289859 654804 289925 654805
rect 289859 654740 289860 654804
rect 289924 654740 289925 654804
rect 289859 654739 289925 654740
rect 299243 654804 299309 654805
rect 299243 654740 299244 654804
rect 299308 654740 299309 654804
rect 299243 654739 299309 654740
rect 299611 654804 299677 654805
rect 299611 654740 299612 654804
rect 299676 654740 299677 654804
rect 299611 654739 299677 654740
rect 308995 654804 309061 654805
rect 308995 654740 308996 654804
rect 309060 654740 309061 654804
rect 308995 654739 309061 654740
rect 309179 654804 309245 654805
rect 309179 654740 309180 654804
rect 309244 654740 309245 654804
rect 309179 654739 309245 654740
rect 318563 654804 318629 654805
rect 318563 654740 318564 654804
rect 318628 654740 318629 654804
rect 318563 654739 318629 654740
rect 318931 654804 318997 654805
rect 318931 654740 318932 654804
rect 318996 654740 318997 654804
rect 318931 654739 318997 654740
rect 328315 654804 328381 654805
rect 328315 654740 328316 654804
rect 328380 654740 328381 654804
rect 328315 654739 328381 654740
rect 328499 654804 328565 654805
rect 328499 654740 328500 654804
rect 328564 654740 328565 654804
rect 328499 654739 328565 654740
rect 337883 654804 337949 654805
rect 337883 654740 337884 654804
rect 337948 654740 337949 654804
rect 337883 654739 337949 654740
rect 338251 654804 338317 654805
rect 338251 654740 338252 654804
rect 338316 654740 338317 654804
rect 338251 654739 338317 654740
rect 347635 654804 347701 654805
rect 347635 654740 347636 654804
rect 347700 654740 347701 654804
rect 347635 654739 347701 654740
rect 347819 654804 347885 654805
rect 347819 654740 347820 654804
rect 347884 654740 347885 654804
rect 347819 654739 347885 654740
rect 357203 654804 357269 654805
rect 357203 654740 357204 654804
rect 357268 654740 357269 654804
rect 357203 654739 357269 654740
rect 357571 654804 357637 654805
rect 357571 654740 357572 654804
rect 357636 654740 357637 654804
rect 357571 654739 357637 654740
rect 366955 654804 367021 654805
rect 366955 654740 366956 654804
rect 367020 654740 367021 654804
rect 366955 654739 367021 654740
rect 367139 654804 367205 654805
rect 367139 654740 367140 654804
rect 367204 654740 367205 654804
rect 367139 654739 367205 654740
rect 376523 654804 376589 654805
rect 376523 654740 376524 654804
rect 376588 654740 376589 654804
rect 376523 654739 376589 654740
rect 222334 653309 222394 654739
rect 231718 654150 231778 654739
rect 231902 654150 231962 654739
rect 231718 654090 231962 654150
rect 241286 654150 241346 654739
rect 241654 654150 241714 654739
rect 241286 654090 241714 654150
rect 251038 654150 251098 654739
rect 251222 654150 251282 654739
rect 251038 654090 251282 654150
rect 260606 654150 260666 654739
rect 260974 654150 261034 654739
rect 260606 654090 261034 654150
rect 270358 654150 270418 654739
rect 270542 654150 270602 654739
rect 270358 654090 270602 654150
rect 279926 654150 279986 654739
rect 280294 654150 280354 654739
rect 279926 654090 280354 654150
rect 289678 654150 289738 654739
rect 289862 654150 289922 654739
rect 289678 654090 289922 654150
rect 299246 654150 299306 654739
rect 299614 654150 299674 654739
rect 299246 654090 299674 654150
rect 308998 654150 309058 654739
rect 309182 654150 309242 654739
rect 308998 654090 309242 654150
rect 318566 654150 318626 654739
rect 318934 654150 318994 654739
rect 318566 654090 318994 654150
rect 328318 654150 328378 654739
rect 328502 654150 328562 654739
rect 328318 654090 328562 654150
rect 337886 654150 337946 654739
rect 338254 654150 338314 654739
rect 337886 654090 338314 654150
rect 347638 654150 347698 654739
rect 347822 654150 347882 654739
rect 347638 654090 347882 654150
rect 357206 654150 357266 654739
rect 357574 654150 357634 654739
rect 357206 654090 357634 654150
rect 366958 654150 367018 654739
rect 367142 654150 367202 654739
rect 366958 654090 367202 654150
rect 376526 654150 376586 654739
rect 376894 654150 376954 655011
rect 376526 654090 376954 654150
rect 392166 653989 392226 655011
rect 504406 654397 504466 655011
rect 504403 654396 504469 654397
rect 504403 654332 504404 654396
rect 504468 654332 504469 654396
rect 504403 654331 504469 654332
rect 512134 654261 512194 655011
rect 512131 654260 512197 654261
rect 512131 654196 512132 654260
rect 512196 654196 512197 654260
rect 512131 654195 512197 654196
rect 392163 653988 392229 653989
rect 392163 653924 392164 653988
rect 392228 653924 392229 653988
rect 392163 653923 392229 653924
rect 523542 653717 523602 655011
rect 523539 653716 523605 653717
rect 523539 653652 523540 653716
rect 523604 653652 523605 653716
rect 523539 653651 523605 653652
rect 536790 653581 536850 655011
rect 536787 653580 536853 653581
rect 536787 653516 536788 653580
rect 536852 653516 536853 653580
rect 536787 653515 536853 653516
rect 222331 653308 222397 653309
rect 222331 653244 222332 653308
rect 222396 653244 222397 653308
rect 222331 653243 222397 653244
rect 222515 653308 222581 653309
rect 222515 653244 222516 653308
rect 222580 653244 222581 653308
rect 222515 653243 222581 653244
rect 222518 653170 222578 653243
rect 221966 653110 222578 653170
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 47008 651454 47328 651486
rect 47008 651218 47050 651454
rect 47286 651218 47328 651454
rect 47008 651134 47328 651218
rect 47008 650898 47050 651134
rect 47286 650898 47328 651134
rect 47008 650866 47328 650898
rect 77728 651454 78048 651486
rect 77728 651218 77770 651454
rect 78006 651218 78048 651454
rect 77728 651134 78048 651218
rect 77728 650898 77770 651134
rect 78006 650898 78048 651134
rect 77728 650866 78048 650898
rect 108448 651454 108768 651486
rect 108448 651218 108490 651454
rect 108726 651218 108768 651454
rect 108448 651134 108768 651218
rect 108448 650898 108490 651134
rect 108726 650898 108768 651134
rect 108448 650866 108768 650898
rect 139168 651454 139488 651486
rect 139168 651218 139210 651454
rect 139446 651218 139488 651454
rect 139168 651134 139488 651218
rect 139168 650898 139210 651134
rect 139446 650898 139488 651134
rect 139168 650866 139488 650898
rect 169888 651454 170208 651486
rect 169888 651218 169930 651454
rect 170166 651218 170208 651454
rect 169888 651134 170208 651218
rect 169888 650898 169930 651134
rect 170166 650898 170208 651134
rect 169888 650866 170208 650898
rect 200608 651454 200928 651486
rect 200608 651218 200650 651454
rect 200886 651218 200928 651454
rect 200608 651134 200928 651218
rect 200608 650898 200650 651134
rect 200886 650898 200928 651134
rect 200608 650866 200928 650898
rect 231328 651454 231648 651486
rect 231328 651218 231370 651454
rect 231606 651218 231648 651454
rect 231328 651134 231648 651218
rect 231328 650898 231370 651134
rect 231606 650898 231648 651134
rect 231328 650866 231648 650898
rect 262048 651454 262368 651486
rect 262048 651218 262090 651454
rect 262326 651218 262368 651454
rect 262048 651134 262368 651218
rect 262048 650898 262090 651134
rect 262326 650898 262368 651134
rect 262048 650866 262368 650898
rect 292768 651454 293088 651486
rect 292768 651218 292810 651454
rect 293046 651218 293088 651454
rect 292768 651134 293088 651218
rect 292768 650898 292810 651134
rect 293046 650898 293088 651134
rect 292768 650866 293088 650898
rect 323488 651454 323808 651486
rect 323488 651218 323530 651454
rect 323766 651218 323808 651454
rect 323488 651134 323808 651218
rect 323488 650898 323530 651134
rect 323766 650898 323808 651134
rect 323488 650866 323808 650898
rect 354208 651454 354528 651486
rect 354208 651218 354250 651454
rect 354486 651218 354528 651454
rect 354208 651134 354528 651218
rect 354208 650898 354250 651134
rect 354486 650898 354528 651134
rect 354208 650866 354528 650898
rect 384928 651454 385248 651486
rect 384928 651218 384970 651454
rect 385206 651218 385248 651454
rect 384928 651134 385248 651218
rect 384928 650898 384970 651134
rect 385206 650898 385248 651134
rect 384928 650866 385248 650898
rect 415648 651454 415968 651486
rect 415648 651218 415690 651454
rect 415926 651218 415968 651454
rect 415648 651134 415968 651218
rect 415648 650898 415690 651134
rect 415926 650898 415968 651134
rect 415648 650866 415968 650898
rect 446368 651454 446688 651486
rect 446368 651218 446410 651454
rect 446646 651218 446688 651454
rect 446368 651134 446688 651218
rect 446368 650898 446410 651134
rect 446646 650898 446688 651134
rect 446368 650866 446688 650898
rect 477088 651454 477408 651486
rect 477088 651218 477130 651454
rect 477366 651218 477408 651454
rect 477088 651134 477408 651218
rect 477088 650898 477130 651134
rect 477366 650898 477408 651134
rect 477088 650866 477408 650898
rect 507808 651454 508128 651486
rect 507808 651218 507850 651454
rect 508086 651218 508128 651454
rect 507808 651134 508128 651218
rect 507808 650898 507850 651134
rect 508086 650898 508128 651134
rect 507808 650866 508128 650898
rect 538528 651454 538848 651486
rect 538528 651218 538570 651454
rect 538806 651218 538848 651454
rect 538528 651134 538848 651218
rect 538528 650898 538570 651134
rect 538806 650898 538848 651134
rect 538528 650866 538848 650898
rect 62368 633454 62688 633486
rect 62368 633218 62410 633454
rect 62646 633218 62688 633454
rect 62368 633134 62688 633218
rect 62368 632898 62410 633134
rect 62646 632898 62688 633134
rect 62368 632866 62688 632898
rect 93088 633454 93408 633486
rect 93088 633218 93130 633454
rect 93366 633218 93408 633454
rect 93088 633134 93408 633218
rect 93088 632898 93130 633134
rect 93366 632898 93408 633134
rect 93088 632866 93408 632898
rect 123808 633454 124128 633486
rect 123808 633218 123850 633454
rect 124086 633218 124128 633454
rect 123808 633134 124128 633218
rect 123808 632898 123850 633134
rect 124086 632898 124128 633134
rect 123808 632866 124128 632898
rect 154528 633454 154848 633486
rect 154528 633218 154570 633454
rect 154806 633218 154848 633454
rect 154528 633134 154848 633218
rect 154528 632898 154570 633134
rect 154806 632898 154848 633134
rect 154528 632866 154848 632898
rect 185248 633454 185568 633486
rect 185248 633218 185290 633454
rect 185526 633218 185568 633454
rect 185248 633134 185568 633218
rect 185248 632898 185290 633134
rect 185526 632898 185568 633134
rect 185248 632866 185568 632898
rect 215968 633454 216288 633486
rect 215968 633218 216010 633454
rect 216246 633218 216288 633454
rect 215968 633134 216288 633218
rect 215968 632898 216010 633134
rect 216246 632898 216288 633134
rect 215968 632866 216288 632898
rect 246688 633454 247008 633486
rect 246688 633218 246730 633454
rect 246966 633218 247008 633454
rect 246688 633134 247008 633218
rect 246688 632898 246730 633134
rect 246966 632898 247008 633134
rect 246688 632866 247008 632898
rect 277408 633454 277728 633486
rect 277408 633218 277450 633454
rect 277686 633218 277728 633454
rect 277408 633134 277728 633218
rect 277408 632898 277450 633134
rect 277686 632898 277728 633134
rect 277408 632866 277728 632898
rect 308128 633454 308448 633486
rect 308128 633218 308170 633454
rect 308406 633218 308448 633454
rect 308128 633134 308448 633218
rect 308128 632898 308170 633134
rect 308406 632898 308448 633134
rect 308128 632866 308448 632898
rect 338848 633454 339168 633486
rect 338848 633218 338890 633454
rect 339126 633218 339168 633454
rect 338848 633134 339168 633218
rect 338848 632898 338890 633134
rect 339126 632898 339168 633134
rect 338848 632866 339168 632898
rect 369568 633454 369888 633486
rect 369568 633218 369610 633454
rect 369846 633218 369888 633454
rect 369568 633134 369888 633218
rect 369568 632898 369610 633134
rect 369846 632898 369888 633134
rect 369568 632866 369888 632898
rect 400288 633454 400608 633486
rect 400288 633218 400330 633454
rect 400566 633218 400608 633454
rect 400288 633134 400608 633218
rect 400288 632898 400330 633134
rect 400566 632898 400608 633134
rect 400288 632866 400608 632898
rect 431008 633454 431328 633486
rect 431008 633218 431050 633454
rect 431286 633218 431328 633454
rect 431008 633134 431328 633218
rect 431008 632898 431050 633134
rect 431286 632898 431328 633134
rect 431008 632866 431328 632898
rect 461728 633454 462048 633486
rect 461728 633218 461770 633454
rect 462006 633218 462048 633454
rect 461728 633134 462048 633218
rect 461728 632898 461770 633134
rect 462006 632898 462048 633134
rect 461728 632866 462048 632898
rect 492448 633454 492768 633486
rect 492448 633218 492490 633454
rect 492726 633218 492768 633454
rect 492448 633134 492768 633218
rect 492448 632898 492490 633134
rect 492726 632898 492768 633134
rect 492448 632866 492768 632898
rect 523168 633454 523488 633486
rect 523168 633218 523210 633454
rect 523446 633218 523488 633454
rect 523168 633134 523488 633218
rect 523168 632898 523210 633134
rect 523446 632898 523488 633134
rect 523168 632866 523488 632898
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 47008 615454 47328 615486
rect 47008 615218 47050 615454
rect 47286 615218 47328 615454
rect 47008 615134 47328 615218
rect 47008 614898 47050 615134
rect 47286 614898 47328 615134
rect 47008 614866 47328 614898
rect 77728 615454 78048 615486
rect 77728 615218 77770 615454
rect 78006 615218 78048 615454
rect 77728 615134 78048 615218
rect 77728 614898 77770 615134
rect 78006 614898 78048 615134
rect 77728 614866 78048 614898
rect 108448 615454 108768 615486
rect 108448 615218 108490 615454
rect 108726 615218 108768 615454
rect 108448 615134 108768 615218
rect 108448 614898 108490 615134
rect 108726 614898 108768 615134
rect 108448 614866 108768 614898
rect 139168 615454 139488 615486
rect 139168 615218 139210 615454
rect 139446 615218 139488 615454
rect 139168 615134 139488 615218
rect 139168 614898 139210 615134
rect 139446 614898 139488 615134
rect 139168 614866 139488 614898
rect 169888 615454 170208 615486
rect 169888 615218 169930 615454
rect 170166 615218 170208 615454
rect 169888 615134 170208 615218
rect 169888 614898 169930 615134
rect 170166 614898 170208 615134
rect 169888 614866 170208 614898
rect 200608 615454 200928 615486
rect 200608 615218 200650 615454
rect 200886 615218 200928 615454
rect 200608 615134 200928 615218
rect 200608 614898 200650 615134
rect 200886 614898 200928 615134
rect 200608 614866 200928 614898
rect 231328 615454 231648 615486
rect 231328 615218 231370 615454
rect 231606 615218 231648 615454
rect 231328 615134 231648 615218
rect 231328 614898 231370 615134
rect 231606 614898 231648 615134
rect 231328 614866 231648 614898
rect 262048 615454 262368 615486
rect 262048 615218 262090 615454
rect 262326 615218 262368 615454
rect 262048 615134 262368 615218
rect 262048 614898 262090 615134
rect 262326 614898 262368 615134
rect 262048 614866 262368 614898
rect 292768 615454 293088 615486
rect 292768 615218 292810 615454
rect 293046 615218 293088 615454
rect 292768 615134 293088 615218
rect 292768 614898 292810 615134
rect 293046 614898 293088 615134
rect 292768 614866 293088 614898
rect 323488 615454 323808 615486
rect 323488 615218 323530 615454
rect 323766 615218 323808 615454
rect 323488 615134 323808 615218
rect 323488 614898 323530 615134
rect 323766 614898 323808 615134
rect 323488 614866 323808 614898
rect 354208 615454 354528 615486
rect 354208 615218 354250 615454
rect 354486 615218 354528 615454
rect 354208 615134 354528 615218
rect 354208 614898 354250 615134
rect 354486 614898 354528 615134
rect 354208 614866 354528 614898
rect 384928 615454 385248 615486
rect 384928 615218 384970 615454
rect 385206 615218 385248 615454
rect 384928 615134 385248 615218
rect 384928 614898 384970 615134
rect 385206 614898 385248 615134
rect 384928 614866 385248 614898
rect 415648 615454 415968 615486
rect 415648 615218 415690 615454
rect 415926 615218 415968 615454
rect 415648 615134 415968 615218
rect 415648 614898 415690 615134
rect 415926 614898 415968 615134
rect 415648 614866 415968 614898
rect 446368 615454 446688 615486
rect 446368 615218 446410 615454
rect 446646 615218 446688 615454
rect 446368 615134 446688 615218
rect 446368 614898 446410 615134
rect 446646 614898 446688 615134
rect 446368 614866 446688 614898
rect 477088 615454 477408 615486
rect 477088 615218 477130 615454
rect 477366 615218 477408 615454
rect 477088 615134 477408 615218
rect 477088 614898 477130 615134
rect 477366 614898 477408 615134
rect 477088 614866 477408 614898
rect 507808 615454 508128 615486
rect 507808 615218 507850 615454
rect 508086 615218 508128 615454
rect 507808 615134 508128 615218
rect 507808 614898 507850 615134
rect 508086 614898 508128 615134
rect 507808 614866 508128 614898
rect 538528 615454 538848 615486
rect 538528 615218 538570 615454
rect 538806 615218 538848 615454
rect 538528 615134 538848 615218
rect 538528 614898 538570 615134
rect 538806 614898 538848 615134
rect 538528 614866 538848 614898
rect 62368 597454 62688 597486
rect 62368 597218 62410 597454
rect 62646 597218 62688 597454
rect 62368 597134 62688 597218
rect 62368 596898 62410 597134
rect 62646 596898 62688 597134
rect 62368 596866 62688 596898
rect 93088 597454 93408 597486
rect 93088 597218 93130 597454
rect 93366 597218 93408 597454
rect 93088 597134 93408 597218
rect 93088 596898 93130 597134
rect 93366 596898 93408 597134
rect 93088 596866 93408 596898
rect 123808 597454 124128 597486
rect 123808 597218 123850 597454
rect 124086 597218 124128 597454
rect 123808 597134 124128 597218
rect 123808 596898 123850 597134
rect 124086 596898 124128 597134
rect 123808 596866 124128 596898
rect 154528 597454 154848 597486
rect 154528 597218 154570 597454
rect 154806 597218 154848 597454
rect 154528 597134 154848 597218
rect 154528 596898 154570 597134
rect 154806 596898 154848 597134
rect 154528 596866 154848 596898
rect 185248 597454 185568 597486
rect 185248 597218 185290 597454
rect 185526 597218 185568 597454
rect 185248 597134 185568 597218
rect 185248 596898 185290 597134
rect 185526 596898 185568 597134
rect 185248 596866 185568 596898
rect 215968 597454 216288 597486
rect 215968 597218 216010 597454
rect 216246 597218 216288 597454
rect 215968 597134 216288 597218
rect 215968 596898 216010 597134
rect 216246 596898 216288 597134
rect 215968 596866 216288 596898
rect 246688 597454 247008 597486
rect 246688 597218 246730 597454
rect 246966 597218 247008 597454
rect 246688 597134 247008 597218
rect 246688 596898 246730 597134
rect 246966 596898 247008 597134
rect 246688 596866 247008 596898
rect 277408 597454 277728 597486
rect 277408 597218 277450 597454
rect 277686 597218 277728 597454
rect 277408 597134 277728 597218
rect 277408 596898 277450 597134
rect 277686 596898 277728 597134
rect 277408 596866 277728 596898
rect 308128 597454 308448 597486
rect 308128 597218 308170 597454
rect 308406 597218 308448 597454
rect 308128 597134 308448 597218
rect 308128 596898 308170 597134
rect 308406 596898 308448 597134
rect 308128 596866 308448 596898
rect 338848 597454 339168 597486
rect 338848 597218 338890 597454
rect 339126 597218 339168 597454
rect 338848 597134 339168 597218
rect 338848 596898 338890 597134
rect 339126 596898 339168 597134
rect 338848 596866 339168 596898
rect 369568 597454 369888 597486
rect 369568 597218 369610 597454
rect 369846 597218 369888 597454
rect 369568 597134 369888 597218
rect 369568 596898 369610 597134
rect 369846 596898 369888 597134
rect 369568 596866 369888 596898
rect 400288 597454 400608 597486
rect 400288 597218 400330 597454
rect 400566 597218 400608 597454
rect 400288 597134 400608 597218
rect 400288 596898 400330 597134
rect 400566 596898 400608 597134
rect 400288 596866 400608 596898
rect 431008 597454 431328 597486
rect 431008 597218 431050 597454
rect 431286 597218 431328 597454
rect 431008 597134 431328 597218
rect 431008 596898 431050 597134
rect 431286 596898 431328 597134
rect 431008 596866 431328 596898
rect 461728 597454 462048 597486
rect 461728 597218 461770 597454
rect 462006 597218 462048 597454
rect 461728 597134 462048 597218
rect 461728 596898 461770 597134
rect 462006 596898 462048 597134
rect 461728 596866 462048 596898
rect 492448 597454 492768 597486
rect 492448 597218 492490 597454
rect 492726 597218 492768 597454
rect 492448 597134 492768 597218
rect 492448 596898 492490 597134
rect 492726 596898 492768 597134
rect 492448 596866 492768 596898
rect 523168 597454 523488 597486
rect 523168 597218 523210 597454
rect 523446 597218 523488 597454
rect 523168 597134 523488 597218
rect 523168 596898 523210 597134
rect 523446 596898 523488 597134
rect 523168 596866 523488 596898
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 47008 579454 47328 579486
rect 47008 579218 47050 579454
rect 47286 579218 47328 579454
rect 47008 579134 47328 579218
rect 47008 578898 47050 579134
rect 47286 578898 47328 579134
rect 47008 578866 47328 578898
rect 77728 579454 78048 579486
rect 77728 579218 77770 579454
rect 78006 579218 78048 579454
rect 77728 579134 78048 579218
rect 77728 578898 77770 579134
rect 78006 578898 78048 579134
rect 77728 578866 78048 578898
rect 108448 579454 108768 579486
rect 108448 579218 108490 579454
rect 108726 579218 108768 579454
rect 108448 579134 108768 579218
rect 108448 578898 108490 579134
rect 108726 578898 108768 579134
rect 108448 578866 108768 578898
rect 139168 579454 139488 579486
rect 139168 579218 139210 579454
rect 139446 579218 139488 579454
rect 139168 579134 139488 579218
rect 139168 578898 139210 579134
rect 139446 578898 139488 579134
rect 139168 578866 139488 578898
rect 169888 579454 170208 579486
rect 169888 579218 169930 579454
rect 170166 579218 170208 579454
rect 169888 579134 170208 579218
rect 169888 578898 169930 579134
rect 170166 578898 170208 579134
rect 169888 578866 170208 578898
rect 200608 579454 200928 579486
rect 200608 579218 200650 579454
rect 200886 579218 200928 579454
rect 200608 579134 200928 579218
rect 200608 578898 200650 579134
rect 200886 578898 200928 579134
rect 200608 578866 200928 578898
rect 231328 579454 231648 579486
rect 231328 579218 231370 579454
rect 231606 579218 231648 579454
rect 231328 579134 231648 579218
rect 231328 578898 231370 579134
rect 231606 578898 231648 579134
rect 231328 578866 231648 578898
rect 262048 579454 262368 579486
rect 262048 579218 262090 579454
rect 262326 579218 262368 579454
rect 262048 579134 262368 579218
rect 262048 578898 262090 579134
rect 262326 578898 262368 579134
rect 262048 578866 262368 578898
rect 292768 579454 293088 579486
rect 292768 579218 292810 579454
rect 293046 579218 293088 579454
rect 292768 579134 293088 579218
rect 292768 578898 292810 579134
rect 293046 578898 293088 579134
rect 292768 578866 293088 578898
rect 323488 579454 323808 579486
rect 323488 579218 323530 579454
rect 323766 579218 323808 579454
rect 323488 579134 323808 579218
rect 323488 578898 323530 579134
rect 323766 578898 323808 579134
rect 323488 578866 323808 578898
rect 354208 579454 354528 579486
rect 354208 579218 354250 579454
rect 354486 579218 354528 579454
rect 354208 579134 354528 579218
rect 354208 578898 354250 579134
rect 354486 578898 354528 579134
rect 354208 578866 354528 578898
rect 384928 579454 385248 579486
rect 384928 579218 384970 579454
rect 385206 579218 385248 579454
rect 384928 579134 385248 579218
rect 384928 578898 384970 579134
rect 385206 578898 385248 579134
rect 384928 578866 385248 578898
rect 415648 579454 415968 579486
rect 415648 579218 415690 579454
rect 415926 579218 415968 579454
rect 415648 579134 415968 579218
rect 415648 578898 415690 579134
rect 415926 578898 415968 579134
rect 415648 578866 415968 578898
rect 446368 579454 446688 579486
rect 446368 579218 446410 579454
rect 446646 579218 446688 579454
rect 446368 579134 446688 579218
rect 446368 578898 446410 579134
rect 446646 578898 446688 579134
rect 446368 578866 446688 578898
rect 477088 579454 477408 579486
rect 477088 579218 477130 579454
rect 477366 579218 477408 579454
rect 477088 579134 477408 579218
rect 477088 578898 477130 579134
rect 477366 578898 477408 579134
rect 477088 578866 477408 578898
rect 507808 579454 508128 579486
rect 507808 579218 507850 579454
rect 508086 579218 508128 579454
rect 507808 579134 508128 579218
rect 507808 578898 507850 579134
rect 508086 578898 508128 579134
rect 507808 578866 508128 578898
rect 538528 579454 538848 579486
rect 538528 579218 538570 579454
rect 538806 579218 538848 579454
rect 538528 579134 538848 579218
rect 538528 578898 538570 579134
rect 538806 578898 538848 579134
rect 538528 578866 538848 578898
rect 62368 561454 62688 561486
rect 62368 561218 62410 561454
rect 62646 561218 62688 561454
rect 62368 561134 62688 561218
rect 62368 560898 62410 561134
rect 62646 560898 62688 561134
rect 62368 560866 62688 560898
rect 93088 561454 93408 561486
rect 93088 561218 93130 561454
rect 93366 561218 93408 561454
rect 93088 561134 93408 561218
rect 93088 560898 93130 561134
rect 93366 560898 93408 561134
rect 93088 560866 93408 560898
rect 123808 561454 124128 561486
rect 123808 561218 123850 561454
rect 124086 561218 124128 561454
rect 123808 561134 124128 561218
rect 123808 560898 123850 561134
rect 124086 560898 124128 561134
rect 123808 560866 124128 560898
rect 154528 561454 154848 561486
rect 154528 561218 154570 561454
rect 154806 561218 154848 561454
rect 154528 561134 154848 561218
rect 154528 560898 154570 561134
rect 154806 560898 154848 561134
rect 154528 560866 154848 560898
rect 185248 561454 185568 561486
rect 185248 561218 185290 561454
rect 185526 561218 185568 561454
rect 185248 561134 185568 561218
rect 185248 560898 185290 561134
rect 185526 560898 185568 561134
rect 185248 560866 185568 560898
rect 215968 561454 216288 561486
rect 215968 561218 216010 561454
rect 216246 561218 216288 561454
rect 215968 561134 216288 561218
rect 215968 560898 216010 561134
rect 216246 560898 216288 561134
rect 215968 560866 216288 560898
rect 246688 561454 247008 561486
rect 246688 561218 246730 561454
rect 246966 561218 247008 561454
rect 246688 561134 247008 561218
rect 246688 560898 246730 561134
rect 246966 560898 247008 561134
rect 246688 560866 247008 560898
rect 277408 561454 277728 561486
rect 277408 561218 277450 561454
rect 277686 561218 277728 561454
rect 277408 561134 277728 561218
rect 277408 560898 277450 561134
rect 277686 560898 277728 561134
rect 277408 560866 277728 560898
rect 308128 561454 308448 561486
rect 308128 561218 308170 561454
rect 308406 561218 308448 561454
rect 308128 561134 308448 561218
rect 308128 560898 308170 561134
rect 308406 560898 308448 561134
rect 308128 560866 308448 560898
rect 338848 561454 339168 561486
rect 338848 561218 338890 561454
rect 339126 561218 339168 561454
rect 338848 561134 339168 561218
rect 338848 560898 338890 561134
rect 339126 560898 339168 561134
rect 338848 560866 339168 560898
rect 369568 561454 369888 561486
rect 369568 561218 369610 561454
rect 369846 561218 369888 561454
rect 369568 561134 369888 561218
rect 369568 560898 369610 561134
rect 369846 560898 369888 561134
rect 369568 560866 369888 560898
rect 400288 561454 400608 561486
rect 400288 561218 400330 561454
rect 400566 561218 400608 561454
rect 400288 561134 400608 561218
rect 400288 560898 400330 561134
rect 400566 560898 400608 561134
rect 400288 560866 400608 560898
rect 431008 561454 431328 561486
rect 431008 561218 431050 561454
rect 431286 561218 431328 561454
rect 431008 561134 431328 561218
rect 431008 560898 431050 561134
rect 431286 560898 431328 561134
rect 431008 560866 431328 560898
rect 461728 561454 462048 561486
rect 461728 561218 461770 561454
rect 462006 561218 462048 561454
rect 461728 561134 462048 561218
rect 461728 560898 461770 561134
rect 462006 560898 462048 561134
rect 461728 560866 462048 560898
rect 492448 561454 492768 561486
rect 492448 561218 492490 561454
rect 492726 561218 492768 561454
rect 492448 561134 492768 561218
rect 492448 560898 492490 561134
rect 492726 560898 492768 561134
rect 492448 560866 492768 560898
rect 523168 561454 523488 561486
rect 523168 561218 523210 561454
rect 523446 561218 523488 561454
rect 523168 561134 523488 561218
rect 523168 560898 523210 561134
rect 523446 560898 523488 561134
rect 523168 560866 523488 560898
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 47008 543454 47328 543486
rect 47008 543218 47050 543454
rect 47286 543218 47328 543454
rect 47008 543134 47328 543218
rect 47008 542898 47050 543134
rect 47286 542898 47328 543134
rect 47008 542866 47328 542898
rect 77728 543454 78048 543486
rect 77728 543218 77770 543454
rect 78006 543218 78048 543454
rect 77728 543134 78048 543218
rect 77728 542898 77770 543134
rect 78006 542898 78048 543134
rect 77728 542866 78048 542898
rect 108448 543454 108768 543486
rect 108448 543218 108490 543454
rect 108726 543218 108768 543454
rect 108448 543134 108768 543218
rect 108448 542898 108490 543134
rect 108726 542898 108768 543134
rect 108448 542866 108768 542898
rect 139168 543454 139488 543486
rect 139168 543218 139210 543454
rect 139446 543218 139488 543454
rect 139168 543134 139488 543218
rect 139168 542898 139210 543134
rect 139446 542898 139488 543134
rect 139168 542866 139488 542898
rect 169888 543454 170208 543486
rect 169888 543218 169930 543454
rect 170166 543218 170208 543454
rect 169888 543134 170208 543218
rect 169888 542898 169930 543134
rect 170166 542898 170208 543134
rect 169888 542866 170208 542898
rect 200608 543454 200928 543486
rect 200608 543218 200650 543454
rect 200886 543218 200928 543454
rect 200608 543134 200928 543218
rect 200608 542898 200650 543134
rect 200886 542898 200928 543134
rect 200608 542866 200928 542898
rect 231328 543454 231648 543486
rect 231328 543218 231370 543454
rect 231606 543218 231648 543454
rect 231328 543134 231648 543218
rect 231328 542898 231370 543134
rect 231606 542898 231648 543134
rect 231328 542866 231648 542898
rect 262048 543454 262368 543486
rect 262048 543218 262090 543454
rect 262326 543218 262368 543454
rect 262048 543134 262368 543218
rect 262048 542898 262090 543134
rect 262326 542898 262368 543134
rect 262048 542866 262368 542898
rect 292768 543454 293088 543486
rect 292768 543218 292810 543454
rect 293046 543218 293088 543454
rect 292768 543134 293088 543218
rect 292768 542898 292810 543134
rect 293046 542898 293088 543134
rect 292768 542866 293088 542898
rect 323488 543454 323808 543486
rect 323488 543218 323530 543454
rect 323766 543218 323808 543454
rect 323488 543134 323808 543218
rect 323488 542898 323530 543134
rect 323766 542898 323808 543134
rect 323488 542866 323808 542898
rect 354208 543454 354528 543486
rect 354208 543218 354250 543454
rect 354486 543218 354528 543454
rect 354208 543134 354528 543218
rect 354208 542898 354250 543134
rect 354486 542898 354528 543134
rect 354208 542866 354528 542898
rect 384928 543454 385248 543486
rect 384928 543218 384970 543454
rect 385206 543218 385248 543454
rect 384928 543134 385248 543218
rect 384928 542898 384970 543134
rect 385206 542898 385248 543134
rect 384928 542866 385248 542898
rect 415648 543454 415968 543486
rect 415648 543218 415690 543454
rect 415926 543218 415968 543454
rect 415648 543134 415968 543218
rect 415648 542898 415690 543134
rect 415926 542898 415968 543134
rect 415648 542866 415968 542898
rect 446368 543454 446688 543486
rect 446368 543218 446410 543454
rect 446646 543218 446688 543454
rect 446368 543134 446688 543218
rect 446368 542898 446410 543134
rect 446646 542898 446688 543134
rect 446368 542866 446688 542898
rect 477088 543454 477408 543486
rect 477088 543218 477130 543454
rect 477366 543218 477408 543454
rect 477088 543134 477408 543218
rect 477088 542898 477130 543134
rect 477366 542898 477408 543134
rect 477088 542866 477408 542898
rect 507808 543454 508128 543486
rect 507808 543218 507850 543454
rect 508086 543218 508128 543454
rect 507808 543134 508128 543218
rect 507808 542898 507850 543134
rect 508086 542898 508128 543134
rect 507808 542866 508128 542898
rect 538528 543454 538848 543486
rect 538528 543218 538570 543454
rect 538806 543218 538848 543454
rect 538528 543134 538848 543218
rect 538528 542898 538570 543134
rect 538806 542898 538848 543134
rect 538528 542866 538848 542898
rect 62368 525454 62688 525486
rect 62368 525218 62410 525454
rect 62646 525218 62688 525454
rect 62368 525134 62688 525218
rect 62368 524898 62410 525134
rect 62646 524898 62688 525134
rect 62368 524866 62688 524898
rect 93088 525454 93408 525486
rect 93088 525218 93130 525454
rect 93366 525218 93408 525454
rect 93088 525134 93408 525218
rect 93088 524898 93130 525134
rect 93366 524898 93408 525134
rect 93088 524866 93408 524898
rect 123808 525454 124128 525486
rect 123808 525218 123850 525454
rect 124086 525218 124128 525454
rect 123808 525134 124128 525218
rect 123808 524898 123850 525134
rect 124086 524898 124128 525134
rect 123808 524866 124128 524898
rect 154528 525454 154848 525486
rect 154528 525218 154570 525454
rect 154806 525218 154848 525454
rect 154528 525134 154848 525218
rect 154528 524898 154570 525134
rect 154806 524898 154848 525134
rect 154528 524866 154848 524898
rect 185248 525454 185568 525486
rect 185248 525218 185290 525454
rect 185526 525218 185568 525454
rect 185248 525134 185568 525218
rect 185248 524898 185290 525134
rect 185526 524898 185568 525134
rect 185248 524866 185568 524898
rect 215968 525454 216288 525486
rect 215968 525218 216010 525454
rect 216246 525218 216288 525454
rect 215968 525134 216288 525218
rect 215968 524898 216010 525134
rect 216246 524898 216288 525134
rect 215968 524866 216288 524898
rect 246688 525454 247008 525486
rect 246688 525218 246730 525454
rect 246966 525218 247008 525454
rect 246688 525134 247008 525218
rect 246688 524898 246730 525134
rect 246966 524898 247008 525134
rect 246688 524866 247008 524898
rect 277408 525454 277728 525486
rect 277408 525218 277450 525454
rect 277686 525218 277728 525454
rect 277408 525134 277728 525218
rect 277408 524898 277450 525134
rect 277686 524898 277728 525134
rect 277408 524866 277728 524898
rect 308128 525454 308448 525486
rect 308128 525218 308170 525454
rect 308406 525218 308448 525454
rect 308128 525134 308448 525218
rect 308128 524898 308170 525134
rect 308406 524898 308448 525134
rect 308128 524866 308448 524898
rect 338848 525454 339168 525486
rect 338848 525218 338890 525454
rect 339126 525218 339168 525454
rect 338848 525134 339168 525218
rect 338848 524898 338890 525134
rect 339126 524898 339168 525134
rect 338848 524866 339168 524898
rect 369568 525454 369888 525486
rect 369568 525218 369610 525454
rect 369846 525218 369888 525454
rect 369568 525134 369888 525218
rect 369568 524898 369610 525134
rect 369846 524898 369888 525134
rect 369568 524866 369888 524898
rect 400288 525454 400608 525486
rect 400288 525218 400330 525454
rect 400566 525218 400608 525454
rect 400288 525134 400608 525218
rect 400288 524898 400330 525134
rect 400566 524898 400608 525134
rect 400288 524866 400608 524898
rect 431008 525454 431328 525486
rect 431008 525218 431050 525454
rect 431286 525218 431328 525454
rect 431008 525134 431328 525218
rect 431008 524898 431050 525134
rect 431286 524898 431328 525134
rect 431008 524866 431328 524898
rect 461728 525454 462048 525486
rect 461728 525218 461770 525454
rect 462006 525218 462048 525454
rect 461728 525134 462048 525218
rect 461728 524898 461770 525134
rect 462006 524898 462048 525134
rect 461728 524866 462048 524898
rect 492448 525454 492768 525486
rect 492448 525218 492490 525454
rect 492726 525218 492768 525454
rect 492448 525134 492768 525218
rect 492448 524898 492490 525134
rect 492726 524898 492768 525134
rect 492448 524866 492768 524898
rect 523168 525454 523488 525486
rect 523168 525218 523210 525454
rect 523446 525218 523488 525454
rect 523168 525134 523488 525218
rect 523168 524898 523210 525134
rect 523446 524898 523488 525134
rect 523168 524866 523488 524898
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 47008 507454 47328 507486
rect 47008 507218 47050 507454
rect 47286 507218 47328 507454
rect 47008 507134 47328 507218
rect 47008 506898 47050 507134
rect 47286 506898 47328 507134
rect 47008 506866 47328 506898
rect 77728 507454 78048 507486
rect 77728 507218 77770 507454
rect 78006 507218 78048 507454
rect 77728 507134 78048 507218
rect 77728 506898 77770 507134
rect 78006 506898 78048 507134
rect 77728 506866 78048 506898
rect 108448 507454 108768 507486
rect 108448 507218 108490 507454
rect 108726 507218 108768 507454
rect 108448 507134 108768 507218
rect 108448 506898 108490 507134
rect 108726 506898 108768 507134
rect 108448 506866 108768 506898
rect 139168 507454 139488 507486
rect 139168 507218 139210 507454
rect 139446 507218 139488 507454
rect 139168 507134 139488 507218
rect 139168 506898 139210 507134
rect 139446 506898 139488 507134
rect 139168 506866 139488 506898
rect 169888 507454 170208 507486
rect 169888 507218 169930 507454
rect 170166 507218 170208 507454
rect 169888 507134 170208 507218
rect 169888 506898 169930 507134
rect 170166 506898 170208 507134
rect 169888 506866 170208 506898
rect 200608 507454 200928 507486
rect 200608 507218 200650 507454
rect 200886 507218 200928 507454
rect 200608 507134 200928 507218
rect 200608 506898 200650 507134
rect 200886 506898 200928 507134
rect 200608 506866 200928 506898
rect 231328 507454 231648 507486
rect 231328 507218 231370 507454
rect 231606 507218 231648 507454
rect 231328 507134 231648 507218
rect 231328 506898 231370 507134
rect 231606 506898 231648 507134
rect 231328 506866 231648 506898
rect 262048 507454 262368 507486
rect 262048 507218 262090 507454
rect 262326 507218 262368 507454
rect 262048 507134 262368 507218
rect 262048 506898 262090 507134
rect 262326 506898 262368 507134
rect 262048 506866 262368 506898
rect 292768 507454 293088 507486
rect 292768 507218 292810 507454
rect 293046 507218 293088 507454
rect 292768 507134 293088 507218
rect 292768 506898 292810 507134
rect 293046 506898 293088 507134
rect 292768 506866 293088 506898
rect 323488 507454 323808 507486
rect 323488 507218 323530 507454
rect 323766 507218 323808 507454
rect 323488 507134 323808 507218
rect 323488 506898 323530 507134
rect 323766 506898 323808 507134
rect 323488 506866 323808 506898
rect 354208 507454 354528 507486
rect 354208 507218 354250 507454
rect 354486 507218 354528 507454
rect 354208 507134 354528 507218
rect 354208 506898 354250 507134
rect 354486 506898 354528 507134
rect 354208 506866 354528 506898
rect 384928 507454 385248 507486
rect 384928 507218 384970 507454
rect 385206 507218 385248 507454
rect 384928 507134 385248 507218
rect 384928 506898 384970 507134
rect 385206 506898 385248 507134
rect 384928 506866 385248 506898
rect 415648 507454 415968 507486
rect 415648 507218 415690 507454
rect 415926 507218 415968 507454
rect 415648 507134 415968 507218
rect 415648 506898 415690 507134
rect 415926 506898 415968 507134
rect 415648 506866 415968 506898
rect 446368 507454 446688 507486
rect 446368 507218 446410 507454
rect 446646 507218 446688 507454
rect 446368 507134 446688 507218
rect 446368 506898 446410 507134
rect 446646 506898 446688 507134
rect 446368 506866 446688 506898
rect 477088 507454 477408 507486
rect 477088 507218 477130 507454
rect 477366 507218 477408 507454
rect 477088 507134 477408 507218
rect 477088 506898 477130 507134
rect 477366 506898 477408 507134
rect 477088 506866 477408 506898
rect 507808 507454 508128 507486
rect 507808 507218 507850 507454
rect 508086 507218 508128 507454
rect 507808 507134 508128 507218
rect 507808 506898 507850 507134
rect 508086 506898 508128 507134
rect 507808 506866 508128 506898
rect 538528 507454 538848 507486
rect 538528 507218 538570 507454
rect 538806 507218 538848 507454
rect 538528 507134 538848 507218
rect 538528 506898 538570 507134
rect 538806 506898 538848 507134
rect 538528 506866 538848 506898
rect 62368 489454 62688 489486
rect 62368 489218 62410 489454
rect 62646 489218 62688 489454
rect 62368 489134 62688 489218
rect 62368 488898 62410 489134
rect 62646 488898 62688 489134
rect 62368 488866 62688 488898
rect 93088 489454 93408 489486
rect 93088 489218 93130 489454
rect 93366 489218 93408 489454
rect 93088 489134 93408 489218
rect 93088 488898 93130 489134
rect 93366 488898 93408 489134
rect 93088 488866 93408 488898
rect 123808 489454 124128 489486
rect 123808 489218 123850 489454
rect 124086 489218 124128 489454
rect 123808 489134 124128 489218
rect 123808 488898 123850 489134
rect 124086 488898 124128 489134
rect 123808 488866 124128 488898
rect 154528 489454 154848 489486
rect 154528 489218 154570 489454
rect 154806 489218 154848 489454
rect 154528 489134 154848 489218
rect 154528 488898 154570 489134
rect 154806 488898 154848 489134
rect 154528 488866 154848 488898
rect 185248 489454 185568 489486
rect 185248 489218 185290 489454
rect 185526 489218 185568 489454
rect 185248 489134 185568 489218
rect 185248 488898 185290 489134
rect 185526 488898 185568 489134
rect 185248 488866 185568 488898
rect 215968 489454 216288 489486
rect 215968 489218 216010 489454
rect 216246 489218 216288 489454
rect 215968 489134 216288 489218
rect 215968 488898 216010 489134
rect 216246 488898 216288 489134
rect 215968 488866 216288 488898
rect 246688 489454 247008 489486
rect 246688 489218 246730 489454
rect 246966 489218 247008 489454
rect 246688 489134 247008 489218
rect 246688 488898 246730 489134
rect 246966 488898 247008 489134
rect 246688 488866 247008 488898
rect 277408 489454 277728 489486
rect 277408 489218 277450 489454
rect 277686 489218 277728 489454
rect 277408 489134 277728 489218
rect 277408 488898 277450 489134
rect 277686 488898 277728 489134
rect 277408 488866 277728 488898
rect 308128 489454 308448 489486
rect 308128 489218 308170 489454
rect 308406 489218 308448 489454
rect 308128 489134 308448 489218
rect 308128 488898 308170 489134
rect 308406 488898 308448 489134
rect 308128 488866 308448 488898
rect 338848 489454 339168 489486
rect 338848 489218 338890 489454
rect 339126 489218 339168 489454
rect 338848 489134 339168 489218
rect 338848 488898 338890 489134
rect 339126 488898 339168 489134
rect 338848 488866 339168 488898
rect 369568 489454 369888 489486
rect 369568 489218 369610 489454
rect 369846 489218 369888 489454
rect 369568 489134 369888 489218
rect 369568 488898 369610 489134
rect 369846 488898 369888 489134
rect 369568 488866 369888 488898
rect 400288 489454 400608 489486
rect 400288 489218 400330 489454
rect 400566 489218 400608 489454
rect 400288 489134 400608 489218
rect 400288 488898 400330 489134
rect 400566 488898 400608 489134
rect 400288 488866 400608 488898
rect 431008 489454 431328 489486
rect 431008 489218 431050 489454
rect 431286 489218 431328 489454
rect 431008 489134 431328 489218
rect 431008 488898 431050 489134
rect 431286 488898 431328 489134
rect 431008 488866 431328 488898
rect 461728 489454 462048 489486
rect 461728 489218 461770 489454
rect 462006 489218 462048 489454
rect 461728 489134 462048 489218
rect 461728 488898 461770 489134
rect 462006 488898 462048 489134
rect 461728 488866 462048 488898
rect 492448 489454 492768 489486
rect 492448 489218 492490 489454
rect 492726 489218 492768 489454
rect 492448 489134 492768 489218
rect 492448 488898 492490 489134
rect 492726 488898 492768 489134
rect 492448 488866 492768 488898
rect 523168 489454 523488 489486
rect 523168 489218 523210 489454
rect 523446 489218 523488 489454
rect 523168 489134 523488 489218
rect 523168 488898 523210 489134
rect 523446 488898 523488 489134
rect 523168 488866 523488 488898
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 47008 471454 47328 471486
rect 47008 471218 47050 471454
rect 47286 471218 47328 471454
rect 47008 471134 47328 471218
rect 47008 470898 47050 471134
rect 47286 470898 47328 471134
rect 47008 470866 47328 470898
rect 77728 471454 78048 471486
rect 77728 471218 77770 471454
rect 78006 471218 78048 471454
rect 77728 471134 78048 471218
rect 77728 470898 77770 471134
rect 78006 470898 78048 471134
rect 77728 470866 78048 470898
rect 108448 471454 108768 471486
rect 108448 471218 108490 471454
rect 108726 471218 108768 471454
rect 108448 471134 108768 471218
rect 108448 470898 108490 471134
rect 108726 470898 108768 471134
rect 108448 470866 108768 470898
rect 139168 471454 139488 471486
rect 139168 471218 139210 471454
rect 139446 471218 139488 471454
rect 139168 471134 139488 471218
rect 139168 470898 139210 471134
rect 139446 470898 139488 471134
rect 139168 470866 139488 470898
rect 169888 471454 170208 471486
rect 169888 471218 169930 471454
rect 170166 471218 170208 471454
rect 169888 471134 170208 471218
rect 169888 470898 169930 471134
rect 170166 470898 170208 471134
rect 169888 470866 170208 470898
rect 200608 471454 200928 471486
rect 200608 471218 200650 471454
rect 200886 471218 200928 471454
rect 200608 471134 200928 471218
rect 200608 470898 200650 471134
rect 200886 470898 200928 471134
rect 200608 470866 200928 470898
rect 231328 471454 231648 471486
rect 231328 471218 231370 471454
rect 231606 471218 231648 471454
rect 231328 471134 231648 471218
rect 231328 470898 231370 471134
rect 231606 470898 231648 471134
rect 231328 470866 231648 470898
rect 262048 471454 262368 471486
rect 262048 471218 262090 471454
rect 262326 471218 262368 471454
rect 262048 471134 262368 471218
rect 262048 470898 262090 471134
rect 262326 470898 262368 471134
rect 262048 470866 262368 470898
rect 292768 471454 293088 471486
rect 292768 471218 292810 471454
rect 293046 471218 293088 471454
rect 292768 471134 293088 471218
rect 292768 470898 292810 471134
rect 293046 470898 293088 471134
rect 292768 470866 293088 470898
rect 323488 471454 323808 471486
rect 323488 471218 323530 471454
rect 323766 471218 323808 471454
rect 323488 471134 323808 471218
rect 323488 470898 323530 471134
rect 323766 470898 323808 471134
rect 323488 470866 323808 470898
rect 354208 471454 354528 471486
rect 354208 471218 354250 471454
rect 354486 471218 354528 471454
rect 354208 471134 354528 471218
rect 354208 470898 354250 471134
rect 354486 470898 354528 471134
rect 354208 470866 354528 470898
rect 384928 471454 385248 471486
rect 384928 471218 384970 471454
rect 385206 471218 385248 471454
rect 384928 471134 385248 471218
rect 384928 470898 384970 471134
rect 385206 470898 385248 471134
rect 384928 470866 385248 470898
rect 415648 471454 415968 471486
rect 415648 471218 415690 471454
rect 415926 471218 415968 471454
rect 415648 471134 415968 471218
rect 415648 470898 415690 471134
rect 415926 470898 415968 471134
rect 415648 470866 415968 470898
rect 446368 471454 446688 471486
rect 446368 471218 446410 471454
rect 446646 471218 446688 471454
rect 446368 471134 446688 471218
rect 446368 470898 446410 471134
rect 446646 470898 446688 471134
rect 446368 470866 446688 470898
rect 477088 471454 477408 471486
rect 477088 471218 477130 471454
rect 477366 471218 477408 471454
rect 477088 471134 477408 471218
rect 477088 470898 477130 471134
rect 477366 470898 477408 471134
rect 477088 470866 477408 470898
rect 507808 471454 508128 471486
rect 507808 471218 507850 471454
rect 508086 471218 508128 471454
rect 507808 471134 508128 471218
rect 507808 470898 507850 471134
rect 508086 470898 508128 471134
rect 507808 470866 508128 470898
rect 538528 471454 538848 471486
rect 538528 471218 538570 471454
rect 538806 471218 538848 471454
rect 538528 471134 538848 471218
rect 538528 470898 538570 471134
rect 538806 470898 538848 471134
rect 538528 470866 538848 470898
rect 62368 453454 62688 453486
rect 62368 453218 62410 453454
rect 62646 453218 62688 453454
rect 62368 453134 62688 453218
rect 62368 452898 62410 453134
rect 62646 452898 62688 453134
rect 62368 452866 62688 452898
rect 93088 453454 93408 453486
rect 93088 453218 93130 453454
rect 93366 453218 93408 453454
rect 93088 453134 93408 453218
rect 93088 452898 93130 453134
rect 93366 452898 93408 453134
rect 93088 452866 93408 452898
rect 123808 453454 124128 453486
rect 123808 453218 123850 453454
rect 124086 453218 124128 453454
rect 123808 453134 124128 453218
rect 123808 452898 123850 453134
rect 124086 452898 124128 453134
rect 123808 452866 124128 452898
rect 154528 453454 154848 453486
rect 154528 453218 154570 453454
rect 154806 453218 154848 453454
rect 154528 453134 154848 453218
rect 154528 452898 154570 453134
rect 154806 452898 154848 453134
rect 154528 452866 154848 452898
rect 185248 453454 185568 453486
rect 185248 453218 185290 453454
rect 185526 453218 185568 453454
rect 185248 453134 185568 453218
rect 185248 452898 185290 453134
rect 185526 452898 185568 453134
rect 185248 452866 185568 452898
rect 215968 453454 216288 453486
rect 215968 453218 216010 453454
rect 216246 453218 216288 453454
rect 215968 453134 216288 453218
rect 215968 452898 216010 453134
rect 216246 452898 216288 453134
rect 215968 452866 216288 452898
rect 246688 453454 247008 453486
rect 246688 453218 246730 453454
rect 246966 453218 247008 453454
rect 246688 453134 247008 453218
rect 246688 452898 246730 453134
rect 246966 452898 247008 453134
rect 246688 452866 247008 452898
rect 277408 453454 277728 453486
rect 277408 453218 277450 453454
rect 277686 453218 277728 453454
rect 277408 453134 277728 453218
rect 277408 452898 277450 453134
rect 277686 452898 277728 453134
rect 277408 452866 277728 452898
rect 308128 453454 308448 453486
rect 308128 453218 308170 453454
rect 308406 453218 308448 453454
rect 308128 453134 308448 453218
rect 308128 452898 308170 453134
rect 308406 452898 308448 453134
rect 308128 452866 308448 452898
rect 338848 453454 339168 453486
rect 338848 453218 338890 453454
rect 339126 453218 339168 453454
rect 338848 453134 339168 453218
rect 338848 452898 338890 453134
rect 339126 452898 339168 453134
rect 338848 452866 339168 452898
rect 369568 453454 369888 453486
rect 369568 453218 369610 453454
rect 369846 453218 369888 453454
rect 369568 453134 369888 453218
rect 369568 452898 369610 453134
rect 369846 452898 369888 453134
rect 369568 452866 369888 452898
rect 400288 453454 400608 453486
rect 400288 453218 400330 453454
rect 400566 453218 400608 453454
rect 400288 453134 400608 453218
rect 400288 452898 400330 453134
rect 400566 452898 400608 453134
rect 400288 452866 400608 452898
rect 431008 453454 431328 453486
rect 431008 453218 431050 453454
rect 431286 453218 431328 453454
rect 431008 453134 431328 453218
rect 431008 452898 431050 453134
rect 431286 452898 431328 453134
rect 431008 452866 431328 452898
rect 461728 453454 462048 453486
rect 461728 453218 461770 453454
rect 462006 453218 462048 453454
rect 461728 453134 462048 453218
rect 461728 452898 461770 453134
rect 462006 452898 462048 453134
rect 461728 452866 462048 452898
rect 492448 453454 492768 453486
rect 492448 453218 492490 453454
rect 492726 453218 492768 453454
rect 492448 453134 492768 453218
rect 492448 452898 492490 453134
rect 492726 452898 492768 453134
rect 492448 452866 492768 452898
rect 523168 453454 523488 453486
rect 523168 453218 523210 453454
rect 523446 453218 523488 453454
rect 523168 453134 523488 453218
rect 523168 452898 523210 453134
rect 523446 452898 523488 453134
rect 523168 452866 523488 452898
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 47008 435454 47328 435486
rect 47008 435218 47050 435454
rect 47286 435218 47328 435454
rect 47008 435134 47328 435218
rect 47008 434898 47050 435134
rect 47286 434898 47328 435134
rect 47008 434866 47328 434898
rect 77728 435454 78048 435486
rect 77728 435218 77770 435454
rect 78006 435218 78048 435454
rect 77728 435134 78048 435218
rect 77728 434898 77770 435134
rect 78006 434898 78048 435134
rect 77728 434866 78048 434898
rect 108448 435454 108768 435486
rect 108448 435218 108490 435454
rect 108726 435218 108768 435454
rect 108448 435134 108768 435218
rect 108448 434898 108490 435134
rect 108726 434898 108768 435134
rect 108448 434866 108768 434898
rect 139168 435454 139488 435486
rect 139168 435218 139210 435454
rect 139446 435218 139488 435454
rect 139168 435134 139488 435218
rect 139168 434898 139210 435134
rect 139446 434898 139488 435134
rect 139168 434866 139488 434898
rect 169888 435454 170208 435486
rect 169888 435218 169930 435454
rect 170166 435218 170208 435454
rect 169888 435134 170208 435218
rect 169888 434898 169930 435134
rect 170166 434898 170208 435134
rect 169888 434866 170208 434898
rect 200608 435454 200928 435486
rect 200608 435218 200650 435454
rect 200886 435218 200928 435454
rect 200608 435134 200928 435218
rect 200608 434898 200650 435134
rect 200886 434898 200928 435134
rect 200608 434866 200928 434898
rect 231328 435454 231648 435486
rect 231328 435218 231370 435454
rect 231606 435218 231648 435454
rect 231328 435134 231648 435218
rect 231328 434898 231370 435134
rect 231606 434898 231648 435134
rect 231328 434866 231648 434898
rect 262048 435454 262368 435486
rect 262048 435218 262090 435454
rect 262326 435218 262368 435454
rect 262048 435134 262368 435218
rect 262048 434898 262090 435134
rect 262326 434898 262368 435134
rect 262048 434866 262368 434898
rect 292768 435454 293088 435486
rect 292768 435218 292810 435454
rect 293046 435218 293088 435454
rect 292768 435134 293088 435218
rect 292768 434898 292810 435134
rect 293046 434898 293088 435134
rect 292768 434866 293088 434898
rect 323488 435454 323808 435486
rect 323488 435218 323530 435454
rect 323766 435218 323808 435454
rect 323488 435134 323808 435218
rect 323488 434898 323530 435134
rect 323766 434898 323808 435134
rect 323488 434866 323808 434898
rect 354208 435454 354528 435486
rect 354208 435218 354250 435454
rect 354486 435218 354528 435454
rect 354208 435134 354528 435218
rect 354208 434898 354250 435134
rect 354486 434898 354528 435134
rect 354208 434866 354528 434898
rect 384928 435454 385248 435486
rect 384928 435218 384970 435454
rect 385206 435218 385248 435454
rect 384928 435134 385248 435218
rect 384928 434898 384970 435134
rect 385206 434898 385248 435134
rect 384928 434866 385248 434898
rect 415648 435454 415968 435486
rect 415648 435218 415690 435454
rect 415926 435218 415968 435454
rect 415648 435134 415968 435218
rect 415648 434898 415690 435134
rect 415926 434898 415968 435134
rect 415648 434866 415968 434898
rect 446368 435454 446688 435486
rect 446368 435218 446410 435454
rect 446646 435218 446688 435454
rect 446368 435134 446688 435218
rect 446368 434898 446410 435134
rect 446646 434898 446688 435134
rect 446368 434866 446688 434898
rect 477088 435454 477408 435486
rect 477088 435218 477130 435454
rect 477366 435218 477408 435454
rect 477088 435134 477408 435218
rect 477088 434898 477130 435134
rect 477366 434898 477408 435134
rect 477088 434866 477408 434898
rect 507808 435454 508128 435486
rect 507808 435218 507850 435454
rect 508086 435218 508128 435454
rect 507808 435134 508128 435218
rect 507808 434898 507850 435134
rect 508086 434898 508128 435134
rect 507808 434866 508128 434898
rect 538528 435454 538848 435486
rect 538528 435218 538570 435454
rect 538806 435218 538848 435454
rect 538528 435134 538848 435218
rect 538528 434898 538570 435134
rect 538806 434898 538848 435134
rect 538528 434866 538848 434898
rect 62368 417454 62688 417486
rect 62368 417218 62410 417454
rect 62646 417218 62688 417454
rect 62368 417134 62688 417218
rect 62368 416898 62410 417134
rect 62646 416898 62688 417134
rect 62368 416866 62688 416898
rect 93088 417454 93408 417486
rect 93088 417218 93130 417454
rect 93366 417218 93408 417454
rect 93088 417134 93408 417218
rect 93088 416898 93130 417134
rect 93366 416898 93408 417134
rect 93088 416866 93408 416898
rect 123808 417454 124128 417486
rect 123808 417218 123850 417454
rect 124086 417218 124128 417454
rect 123808 417134 124128 417218
rect 123808 416898 123850 417134
rect 124086 416898 124128 417134
rect 123808 416866 124128 416898
rect 154528 417454 154848 417486
rect 154528 417218 154570 417454
rect 154806 417218 154848 417454
rect 154528 417134 154848 417218
rect 154528 416898 154570 417134
rect 154806 416898 154848 417134
rect 154528 416866 154848 416898
rect 185248 417454 185568 417486
rect 185248 417218 185290 417454
rect 185526 417218 185568 417454
rect 185248 417134 185568 417218
rect 185248 416898 185290 417134
rect 185526 416898 185568 417134
rect 185248 416866 185568 416898
rect 215968 417454 216288 417486
rect 215968 417218 216010 417454
rect 216246 417218 216288 417454
rect 215968 417134 216288 417218
rect 215968 416898 216010 417134
rect 216246 416898 216288 417134
rect 215968 416866 216288 416898
rect 246688 417454 247008 417486
rect 246688 417218 246730 417454
rect 246966 417218 247008 417454
rect 246688 417134 247008 417218
rect 246688 416898 246730 417134
rect 246966 416898 247008 417134
rect 246688 416866 247008 416898
rect 277408 417454 277728 417486
rect 277408 417218 277450 417454
rect 277686 417218 277728 417454
rect 277408 417134 277728 417218
rect 277408 416898 277450 417134
rect 277686 416898 277728 417134
rect 277408 416866 277728 416898
rect 308128 417454 308448 417486
rect 308128 417218 308170 417454
rect 308406 417218 308448 417454
rect 308128 417134 308448 417218
rect 308128 416898 308170 417134
rect 308406 416898 308448 417134
rect 308128 416866 308448 416898
rect 338848 417454 339168 417486
rect 338848 417218 338890 417454
rect 339126 417218 339168 417454
rect 338848 417134 339168 417218
rect 338848 416898 338890 417134
rect 339126 416898 339168 417134
rect 338848 416866 339168 416898
rect 369568 417454 369888 417486
rect 369568 417218 369610 417454
rect 369846 417218 369888 417454
rect 369568 417134 369888 417218
rect 369568 416898 369610 417134
rect 369846 416898 369888 417134
rect 369568 416866 369888 416898
rect 400288 417454 400608 417486
rect 400288 417218 400330 417454
rect 400566 417218 400608 417454
rect 400288 417134 400608 417218
rect 400288 416898 400330 417134
rect 400566 416898 400608 417134
rect 400288 416866 400608 416898
rect 431008 417454 431328 417486
rect 431008 417218 431050 417454
rect 431286 417218 431328 417454
rect 431008 417134 431328 417218
rect 431008 416898 431050 417134
rect 431286 416898 431328 417134
rect 431008 416866 431328 416898
rect 461728 417454 462048 417486
rect 461728 417218 461770 417454
rect 462006 417218 462048 417454
rect 461728 417134 462048 417218
rect 461728 416898 461770 417134
rect 462006 416898 462048 417134
rect 461728 416866 462048 416898
rect 492448 417454 492768 417486
rect 492448 417218 492490 417454
rect 492726 417218 492768 417454
rect 492448 417134 492768 417218
rect 492448 416898 492490 417134
rect 492726 416898 492768 417134
rect 492448 416866 492768 416898
rect 523168 417454 523488 417486
rect 523168 417218 523210 417454
rect 523446 417218 523488 417454
rect 523168 417134 523488 417218
rect 523168 416898 523210 417134
rect 523446 416898 523488 417134
rect 523168 416866 523488 416898
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 47008 399454 47328 399486
rect 47008 399218 47050 399454
rect 47286 399218 47328 399454
rect 47008 399134 47328 399218
rect 47008 398898 47050 399134
rect 47286 398898 47328 399134
rect 47008 398866 47328 398898
rect 77728 399454 78048 399486
rect 77728 399218 77770 399454
rect 78006 399218 78048 399454
rect 77728 399134 78048 399218
rect 77728 398898 77770 399134
rect 78006 398898 78048 399134
rect 77728 398866 78048 398898
rect 108448 399454 108768 399486
rect 108448 399218 108490 399454
rect 108726 399218 108768 399454
rect 108448 399134 108768 399218
rect 108448 398898 108490 399134
rect 108726 398898 108768 399134
rect 108448 398866 108768 398898
rect 139168 399454 139488 399486
rect 139168 399218 139210 399454
rect 139446 399218 139488 399454
rect 139168 399134 139488 399218
rect 139168 398898 139210 399134
rect 139446 398898 139488 399134
rect 139168 398866 139488 398898
rect 169888 399454 170208 399486
rect 169888 399218 169930 399454
rect 170166 399218 170208 399454
rect 169888 399134 170208 399218
rect 169888 398898 169930 399134
rect 170166 398898 170208 399134
rect 169888 398866 170208 398898
rect 200608 399454 200928 399486
rect 200608 399218 200650 399454
rect 200886 399218 200928 399454
rect 200608 399134 200928 399218
rect 200608 398898 200650 399134
rect 200886 398898 200928 399134
rect 200608 398866 200928 398898
rect 231328 399454 231648 399486
rect 231328 399218 231370 399454
rect 231606 399218 231648 399454
rect 231328 399134 231648 399218
rect 231328 398898 231370 399134
rect 231606 398898 231648 399134
rect 231328 398866 231648 398898
rect 262048 399454 262368 399486
rect 262048 399218 262090 399454
rect 262326 399218 262368 399454
rect 262048 399134 262368 399218
rect 262048 398898 262090 399134
rect 262326 398898 262368 399134
rect 262048 398866 262368 398898
rect 292768 399454 293088 399486
rect 292768 399218 292810 399454
rect 293046 399218 293088 399454
rect 292768 399134 293088 399218
rect 292768 398898 292810 399134
rect 293046 398898 293088 399134
rect 292768 398866 293088 398898
rect 323488 399454 323808 399486
rect 323488 399218 323530 399454
rect 323766 399218 323808 399454
rect 323488 399134 323808 399218
rect 323488 398898 323530 399134
rect 323766 398898 323808 399134
rect 323488 398866 323808 398898
rect 354208 399454 354528 399486
rect 354208 399218 354250 399454
rect 354486 399218 354528 399454
rect 354208 399134 354528 399218
rect 354208 398898 354250 399134
rect 354486 398898 354528 399134
rect 354208 398866 354528 398898
rect 384928 399454 385248 399486
rect 384928 399218 384970 399454
rect 385206 399218 385248 399454
rect 384928 399134 385248 399218
rect 384928 398898 384970 399134
rect 385206 398898 385248 399134
rect 384928 398866 385248 398898
rect 415648 399454 415968 399486
rect 415648 399218 415690 399454
rect 415926 399218 415968 399454
rect 415648 399134 415968 399218
rect 415648 398898 415690 399134
rect 415926 398898 415968 399134
rect 415648 398866 415968 398898
rect 446368 399454 446688 399486
rect 446368 399218 446410 399454
rect 446646 399218 446688 399454
rect 446368 399134 446688 399218
rect 446368 398898 446410 399134
rect 446646 398898 446688 399134
rect 446368 398866 446688 398898
rect 477088 399454 477408 399486
rect 477088 399218 477130 399454
rect 477366 399218 477408 399454
rect 477088 399134 477408 399218
rect 477088 398898 477130 399134
rect 477366 398898 477408 399134
rect 477088 398866 477408 398898
rect 507808 399454 508128 399486
rect 507808 399218 507850 399454
rect 508086 399218 508128 399454
rect 507808 399134 508128 399218
rect 507808 398898 507850 399134
rect 508086 398898 508128 399134
rect 507808 398866 508128 398898
rect 538528 399454 538848 399486
rect 538528 399218 538570 399454
rect 538806 399218 538848 399454
rect 538528 399134 538848 399218
rect 538528 398898 538570 399134
rect 538806 398898 538848 399134
rect 538528 398866 538848 398898
rect 62368 381454 62688 381486
rect 62368 381218 62410 381454
rect 62646 381218 62688 381454
rect 62368 381134 62688 381218
rect 62368 380898 62410 381134
rect 62646 380898 62688 381134
rect 62368 380866 62688 380898
rect 93088 381454 93408 381486
rect 93088 381218 93130 381454
rect 93366 381218 93408 381454
rect 93088 381134 93408 381218
rect 93088 380898 93130 381134
rect 93366 380898 93408 381134
rect 93088 380866 93408 380898
rect 123808 381454 124128 381486
rect 123808 381218 123850 381454
rect 124086 381218 124128 381454
rect 123808 381134 124128 381218
rect 123808 380898 123850 381134
rect 124086 380898 124128 381134
rect 123808 380866 124128 380898
rect 154528 381454 154848 381486
rect 154528 381218 154570 381454
rect 154806 381218 154848 381454
rect 154528 381134 154848 381218
rect 154528 380898 154570 381134
rect 154806 380898 154848 381134
rect 154528 380866 154848 380898
rect 185248 381454 185568 381486
rect 185248 381218 185290 381454
rect 185526 381218 185568 381454
rect 185248 381134 185568 381218
rect 185248 380898 185290 381134
rect 185526 380898 185568 381134
rect 185248 380866 185568 380898
rect 215968 381454 216288 381486
rect 215968 381218 216010 381454
rect 216246 381218 216288 381454
rect 215968 381134 216288 381218
rect 215968 380898 216010 381134
rect 216246 380898 216288 381134
rect 215968 380866 216288 380898
rect 246688 381454 247008 381486
rect 246688 381218 246730 381454
rect 246966 381218 247008 381454
rect 246688 381134 247008 381218
rect 246688 380898 246730 381134
rect 246966 380898 247008 381134
rect 246688 380866 247008 380898
rect 277408 381454 277728 381486
rect 277408 381218 277450 381454
rect 277686 381218 277728 381454
rect 277408 381134 277728 381218
rect 277408 380898 277450 381134
rect 277686 380898 277728 381134
rect 277408 380866 277728 380898
rect 308128 381454 308448 381486
rect 308128 381218 308170 381454
rect 308406 381218 308448 381454
rect 308128 381134 308448 381218
rect 308128 380898 308170 381134
rect 308406 380898 308448 381134
rect 308128 380866 308448 380898
rect 338848 381454 339168 381486
rect 338848 381218 338890 381454
rect 339126 381218 339168 381454
rect 338848 381134 339168 381218
rect 338848 380898 338890 381134
rect 339126 380898 339168 381134
rect 338848 380866 339168 380898
rect 369568 381454 369888 381486
rect 369568 381218 369610 381454
rect 369846 381218 369888 381454
rect 369568 381134 369888 381218
rect 369568 380898 369610 381134
rect 369846 380898 369888 381134
rect 369568 380866 369888 380898
rect 400288 381454 400608 381486
rect 400288 381218 400330 381454
rect 400566 381218 400608 381454
rect 400288 381134 400608 381218
rect 400288 380898 400330 381134
rect 400566 380898 400608 381134
rect 400288 380866 400608 380898
rect 431008 381454 431328 381486
rect 431008 381218 431050 381454
rect 431286 381218 431328 381454
rect 431008 381134 431328 381218
rect 431008 380898 431050 381134
rect 431286 380898 431328 381134
rect 431008 380866 431328 380898
rect 461728 381454 462048 381486
rect 461728 381218 461770 381454
rect 462006 381218 462048 381454
rect 461728 381134 462048 381218
rect 461728 380898 461770 381134
rect 462006 380898 462048 381134
rect 461728 380866 462048 380898
rect 492448 381454 492768 381486
rect 492448 381218 492490 381454
rect 492726 381218 492768 381454
rect 492448 381134 492768 381218
rect 492448 380898 492490 381134
rect 492726 380898 492768 381134
rect 492448 380866 492768 380898
rect 523168 381454 523488 381486
rect 523168 381218 523210 381454
rect 523446 381218 523488 381454
rect 523168 381134 523488 381218
rect 523168 380898 523210 381134
rect 523446 380898 523488 381134
rect 523168 380866 523488 380898
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 47008 363454 47328 363486
rect 47008 363218 47050 363454
rect 47286 363218 47328 363454
rect 47008 363134 47328 363218
rect 47008 362898 47050 363134
rect 47286 362898 47328 363134
rect 47008 362866 47328 362898
rect 77728 363454 78048 363486
rect 77728 363218 77770 363454
rect 78006 363218 78048 363454
rect 77728 363134 78048 363218
rect 77728 362898 77770 363134
rect 78006 362898 78048 363134
rect 77728 362866 78048 362898
rect 108448 363454 108768 363486
rect 108448 363218 108490 363454
rect 108726 363218 108768 363454
rect 108448 363134 108768 363218
rect 108448 362898 108490 363134
rect 108726 362898 108768 363134
rect 108448 362866 108768 362898
rect 139168 363454 139488 363486
rect 139168 363218 139210 363454
rect 139446 363218 139488 363454
rect 139168 363134 139488 363218
rect 139168 362898 139210 363134
rect 139446 362898 139488 363134
rect 139168 362866 139488 362898
rect 169888 363454 170208 363486
rect 169888 363218 169930 363454
rect 170166 363218 170208 363454
rect 169888 363134 170208 363218
rect 169888 362898 169930 363134
rect 170166 362898 170208 363134
rect 169888 362866 170208 362898
rect 200608 363454 200928 363486
rect 200608 363218 200650 363454
rect 200886 363218 200928 363454
rect 200608 363134 200928 363218
rect 200608 362898 200650 363134
rect 200886 362898 200928 363134
rect 200608 362866 200928 362898
rect 231328 363454 231648 363486
rect 231328 363218 231370 363454
rect 231606 363218 231648 363454
rect 231328 363134 231648 363218
rect 231328 362898 231370 363134
rect 231606 362898 231648 363134
rect 231328 362866 231648 362898
rect 262048 363454 262368 363486
rect 262048 363218 262090 363454
rect 262326 363218 262368 363454
rect 262048 363134 262368 363218
rect 262048 362898 262090 363134
rect 262326 362898 262368 363134
rect 262048 362866 262368 362898
rect 292768 363454 293088 363486
rect 292768 363218 292810 363454
rect 293046 363218 293088 363454
rect 292768 363134 293088 363218
rect 292768 362898 292810 363134
rect 293046 362898 293088 363134
rect 292768 362866 293088 362898
rect 323488 363454 323808 363486
rect 323488 363218 323530 363454
rect 323766 363218 323808 363454
rect 323488 363134 323808 363218
rect 323488 362898 323530 363134
rect 323766 362898 323808 363134
rect 323488 362866 323808 362898
rect 354208 363454 354528 363486
rect 354208 363218 354250 363454
rect 354486 363218 354528 363454
rect 354208 363134 354528 363218
rect 354208 362898 354250 363134
rect 354486 362898 354528 363134
rect 354208 362866 354528 362898
rect 384928 363454 385248 363486
rect 384928 363218 384970 363454
rect 385206 363218 385248 363454
rect 384928 363134 385248 363218
rect 384928 362898 384970 363134
rect 385206 362898 385248 363134
rect 384928 362866 385248 362898
rect 415648 363454 415968 363486
rect 415648 363218 415690 363454
rect 415926 363218 415968 363454
rect 415648 363134 415968 363218
rect 415648 362898 415690 363134
rect 415926 362898 415968 363134
rect 415648 362866 415968 362898
rect 446368 363454 446688 363486
rect 446368 363218 446410 363454
rect 446646 363218 446688 363454
rect 446368 363134 446688 363218
rect 446368 362898 446410 363134
rect 446646 362898 446688 363134
rect 446368 362866 446688 362898
rect 477088 363454 477408 363486
rect 477088 363218 477130 363454
rect 477366 363218 477408 363454
rect 477088 363134 477408 363218
rect 477088 362898 477130 363134
rect 477366 362898 477408 363134
rect 477088 362866 477408 362898
rect 507808 363454 508128 363486
rect 507808 363218 507850 363454
rect 508086 363218 508128 363454
rect 507808 363134 508128 363218
rect 507808 362898 507850 363134
rect 508086 362898 508128 363134
rect 507808 362866 508128 362898
rect 538528 363454 538848 363486
rect 538528 363218 538570 363454
rect 538806 363218 538848 363454
rect 538528 363134 538848 363218
rect 538528 362898 538570 363134
rect 538806 362898 538848 363134
rect 538528 362866 538848 362898
rect 62368 345454 62688 345486
rect 62368 345218 62410 345454
rect 62646 345218 62688 345454
rect 62368 345134 62688 345218
rect 62368 344898 62410 345134
rect 62646 344898 62688 345134
rect 62368 344866 62688 344898
rect 93088 345454 93408 345486
rect 93088 345218 93130 345454
rect 93366 345218 93408 345454
rect 93088 345134 93408 345218
rect 93088 344898 93130 345134
rect 93366 344898 93408 345134
rect 93088 344866 93408 344898
rect 123808 345454 124128 345486
rect 123808 345218 123850 345454
rect 124086 345218 124128 345454
rect 123808 345134 124128 345218
rect 123808 344898 123850 345134
rect 124086 344898 124128 345134
rect 123808 344866 124128 344898
rect 154528 345454 154848 345486
rect 154528 345218 154570 345454
rect 154806 345218 154848 345454
rect 154528 345134 154848 345218
rect 154528 344898 154570 345134
rect 154806 344898 154848 345134
rect 154528 344866 154848 344898
rect 185248 345454 185568 345486
rect 185248 345218 185290 345454
rect 185526 345218 185568 345454
rect 185248 345134 185568 345218
rect 185248 344898 185290 345134
rect 185526 344898 185568 345134
rect 185248 344866 185568 344898
rect 215968 345454 216288 345486
rect 215968 345218 216010 345454
rect 216246 345218 216288 345454
rect 215968 345134 216288 345218
rect 215968 344898 216010 345134
rect 216246 344898 216288 345134
rect 215968 344866 216288 344898
rect 246688 345454 247008 345486
rect 246688 345218 246730 345454
rect 246966 345218 247008 345454
rect 246688 345134 247008 345218
rect 246688 344898 246730 345134
rect 246966 344898 247008 345134
rect 246688 344866 247008 344898
rect 277408 345454 277728 345486
rect 277408 345218 277450 345454
rect 277686 345218 277728 345454
rect 277408 345134 277728 345218
rect 277408 344898 277450 345134
rect 277686 344898 277728 345134
rect 277408 344866 277728 344898
rect 308128 345454 308448 345486
rect 308128 345218 308170 345454
rect 308406 345218 308448 345454
rect 308128 345134 308448 345218
rect 308128 344898 308170 345134
rect 308406 344898 308448 345134
rect 308128 344866 308448 344898
rect 338848 345454 339168 345486
rect 338848 345218 338890 345454
rect 339126 345218 339168 345454
rect 338848 345134 339168 345218
rect 338848 344898 338890 345134
rect 339126 344898 339168 345134
rect 338848 344866 339168 344898
rect 369568 345454 369888 345486
rect 369568 345218 369610 345454
rect 369846 345218 369888 345454
rect 369568 345134 369888 345218
rect 369568 344898 369610 345134
rect 369846 344898 369888 345134
rect 369568 344866 369888 344898
rect 400288 345454 400608 345486
rect 400288 345218 400330 345454
rect 400566 345218 400608 345454
rect 400288 345134 400608 345218
rect 400288 344898 400330 345134
rect 400566 344898 400608 345134
rect 400288 344866 400608 344898
rect 431008 345454 431328 345486
rect 431008 345218 431050 345454
rect 431286 345218 431328 345454
rect 431008 345134 431328 345218
rect 431008 344898 431050 345134
rect 431286 344898 431328 345134
rect 431008 344866 431328 344898
rect 461728 345454 462048 345486
rect 461728 345218 461770 345454
rect 462006 345218 462048 345454
rect 461728 345134 462048 345218
rect 461728 344898 461770 345134
rect 462006 344898 462048 345134
rect 461728 344866 462048 344898
rect 492448 345454 492768 345486
rect 492448 345218 492490 345454
rect 492726 345218 492768 345454
rect 492448 345134 492768 345218
rect 492448 344898 492490 345134
rect 492726 344898 492768 345134
rect 492448 344866 492768 344898
rect 523168 345454 523488 345486
rect 523168 345218 523210 345454
rect 523446 345218 523488 345454
rect 523168 345134 523488 345218
rect 523168 344898 523210 345134
rect 523446 344898 523488 345134
rect 523168 344866 523488 344898
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 47008 327454 47328 327486
rect 47008 327218 47050 327454
rect 47286 327218 47328 327454
rect 47008 327134 47328 327218
rect 47008 326898 47050 327134
rect 47286 326898 47328 327134
rect 47008 326866 47328 326898
rect 77728 327454 78048 327486
rect 77728 327218 77770 327454
rect 78006 327218 78048 327454
rect 77728 327134 78048 327218
rect 77728 326898 77770 327134
rect 78006 326898 78048 327134
rect 77728 326866 78048 326898
rect 108448 327454 108768 327486
rect 108448 327218 108490 327454
rect 108726 327218 108768 327454
rect 108448 327134 108768 327218
rect 108448 326898 108490 327134
rect 108726 326898 108768 327134
rect 108448 326866 108768 326898
rect 139168 327454 139488 327486
rect 139168 327218 139210 327454
rect 139446 327218 139488 327454
rect 139168 327134 139488 327218
rect 139168 326898 139210 327134
rect 139446 326898 139488 327134
rect 139168 326866 139488 326898
rect 169888 327454 170208 327486
rect 169888 327218 169930 327454
rect 170166 327218 170208 327454
rect 169888 327134 170208 327218
rect 169888 326898 169930 327134
rect 170166 326898 170208 327134
rect 169888 326866 170208 326898
rect 200608 327454 200928 327486
rect 200608 327218 200650 327454
rect 200886 327218 200928 327454
rect 200608 327134 200928 327218
rect 200608 326898 200650 327134
rect 200886 326898 200928 327134
rect 200608 326866 200928 326898
rect 231328 327454 231648 327486
rect 231328 327218 231370 327454
rect 231606 327218 231648 327454
rect 231328 327134 231648 327218
rect 231328 326898 231370 327134
rect 231606 326898 231648 327134
rect 231328 326866 231648 326898
rect 262048 327454 262368 327486
rect 262048 327218 262090 327454
rect 262326 327218 262368 327454
rect 262048 327134 262368 327218
rect 262048 326898 262090 327134
rect 262326 326898 262368 327134
rect 262048 326866 262368 326898
rect 292768 327454 293088 327486
rect 292768 327218 292810 327454
rect 293046 327218 293088 327454
rect 292768 327134 293088 327218
rect 292768 326898 292810 327134
rect 293046 326898 293088 327134
rect 292768 326866 293088 326898
rect 323488 327454 323808 327486
rect 323488 327218 323530 327454
rect 323766 327218 323808 327454
rect 323488 327134 323808 327218
rect 323488 326898 323530 327134
rect 323766 326898 323808 327134
rect 323488 326866 323808 326898
rect 354208 327454 354528 327486
rect 354208 327218 354250 327454
rect 354486 327218 354528 327454
rect 354208 327134 354528 327218
rect 354208 326898 354250 327134
rect 354486 326898 354528 327134
rect 354208 326866 354528 326898
rect 384928 327454 385248 327486
rect 384928 327218 384970 327454
rect 385206 327218 385248 327454
rect 384928 327134 385248 327218
rect 384928 326898 384970 327134
rect 385206 326898 385248 327134
rect 384928 326866 385248 326898
rect 415648 327454 415968 327486
rect 415648 327218 415690 327454
rect 415926 327218 415968 327454
rect 415648 327134 415968 327218
rect 415648 326898 415690 327134
rect 415926 326898 415968 327134
rect 415648 326866 415968 326898
rect 446368 327454 446688 327486
rect 446368 327218 446410 327454
rect 446646 327218 446688 327454
rect 446368 327134 446688 327218
rect 446368 326898 446410 327134
rect 446646 326898 446688 327134
rect 446368 326866 446688 326898
rect 477088 327454 477408 327486
rect 477088 327218 477130 327454
rect 477366 327218 477408 327454
rect 477088 327134 477408 327218
rect 477088 326898 477130 327134
rect 477366 326898 477408 327134
rect 477088 326866 477408 326898
rect 507808 327454 508128 327486
rect 507808 327218 507850 327454
rect 508086 327218 508128 327454
rect 507808 327134 508128 327218
rect 507808 326898 507850 327134
rect 508086 326898 508128 327134
rect 507808 326866 508128 326898
rect 538528 327454 538848 327486
rect 538528 327218 538570 327454
rect 538806 327218 538848 327454
rect 538528 327134 538848 327218
rect 538528 326898 538570 327134
rect 538806 326898 538848 327134
rect 538528 326866 538848 326898
rect 62368 309454 62688 309486
rect 62368 309218 62410 309454
rect 62646 309218 62688 309454
rect 62368 309134 62688 309218
rect 62368 308898 62410 309134
rect 62646 308898 62688 309134
rect 62368 308866 62688 308898
rect 93088 309454 93408 309486
rect 93088 309218 93130 309454
rect 93366 309218 93408 309454
rect 93088 309134 93408 309218
rect 93088 308898 93130 309134
rect 93366 308898 93408 309134
rect 93088 308866 93408 308898
rect 123808 309454 124128 309486
rect 123808 309218 123850 309454
rect 124086 309218 124128 309454
rect 123808 309134 124128 309218
rect 123808 308898 123850 309134
rect 124086 308898 124128 309134
rect 123808 308866 124128 308898
rect 154528 309454 154848 309486
rect 154528 309218 154570 309454
rect 154806 309218 154848 309454
rect 154528 309134 154848 309218
rect 154528 308898 154570 309134
rect 154806 308898 154848 309134
rect 154528 308866 154848 308898
rect 185248 309454 185568 309486
rect 185248 309218 185290 309454
rect 185526 309218 185568 309454
rect 185248 309134 185568 309218
rect 185248 308898 185290 309134
rect 185526 308898 185568 309134
rect 185248 308866 185568 308898
rect 215968 309454 216288 309486
rect 215968 309218 216010 309454
rect 216246 309218 216288 309454
rect 215968 309134 216288 309218
rect 215968 308898 216010 309134
rect 216246 308898 216288 309134
rect 215968 308866 216288 308898
rect 246688 309454 247008 309486
rect 246688 309218 246730 309454
rect 246966 309218 247008 309454
rect 246688 309134 247008 309218
rect 246688 308898 246730 309134
rect 246966 308898 247008 309134
rect 246688 308866 247008 308898
rect 277408 309454 277728 309486
rect 277408 309218 277450 309454
rect 277686 309218 277728 309454
rect 277408 309134 277728 309218
rect 277408 308898 277450 309134
rect 277686 308898 277728 309134
rect 277408 308866 277728 308898
rect 308128 309454 308448 309486
rect 308128 309218 308170 309454
rect 308406 309218 308448 309454
rect 308128 309134 308448 309218
rect 308128 308898 308170 309134
rect 308406 308898 308448 309134
rect 308128 308866 308448 308898
rect 338848 309454 339168 309486
rect 338848 309218 338890 309454
rect 339126 309218 339168 309454
rect 338848 309134 339168 309218
rect 338848 308898 338890 309134
rect 339126 308898 339168 309134
rect 338848 308866 339168 308898
rect 369568 309454 369888 309486
rect 369568 309218 369610 309454
rect 369846 309218 369888 309454
rect 369568 309134 369888 309218
rect 369568 308898 369610 309134
rect 369846 308898 369888 309134
rect 369568 308866 369888 308898
rect 400288 309454 400608 309486
rect 400288 309218 400330 309454
rect 400566 309218 400608 309454
rect 400288 309134 400608 309218
rect 400288 308898 400330 309134
rect 400566 308898 400608 309134
rect 400288 308866 400608 308898
rect 431008 309454 431328 309486
rect 431008 309218 431050 309454
rect 431286 309218 431328 309454
rect 431008 309134 431328 309218
rect 431008 308898 431050 309134
rect 431286 308898 431328 309134
rect 431008 308866 431328 308898
rect 461728 309454 462048 309486
rect 461728 309218 461770 309454
rect 462006 309218 462048 309454
rect 461728 309134 462048 309218
rect 461728 308898 461770 309134
rect 462006 308898 462048 309134
rect 461728 308866 462048 308898
rect 492448 309454 492768 309486
rect 492448 309218 492490 309454
rect 492726 309218 492768 309454
rect 492448 309134 492768 309218
rect 492448 308898 492490 309134
rect 492726 308898 492768 309134
rect 492448 308866 492768 308898
rect 523168 309454 523488 309486
rect 523168 309218 523210 309454
rect 523446 309218 523488 309454
rect 523168 309134 523488 309218
rect 523168 308898 523210 309134
rect 523446 308898 523488 309134
rect 523168 308866 523488 308898
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 47008 291454 47328 291486
rect 47008 291218 47050 291454
rect 47286 291218 47328 291454
rect 47008 291134 47328 291218
rect 47008 290898 47050 291134
rect 47286 290898 47328 291134
rect 47008 290866 47328 290898
rect 77728 291454 78048 291486
rect 77728 291218 77770 291454
rect 78006 291218 78048 291454
rect 77728 291134 78048 291218
rect 77728 290898 77770 291134
rect 78006 290898 78048 291134
rect 77728 290866 78048 290898
rect 108448 291454 108768 291486
rect 108448 291218 108490 291454
rect 108726 291218 108768 291454
rect 108448 291134 108768 291218
rect 108448 290898 108490 291134
rect 108726 290898 108768 291134
rect 108448 290866 108768 290898
rect 139168 291454 139488 291486
rect 139168 291218 139210 291454
rect 139446 291218 139488 291454
rect 139168 291134 139488 291218
rect 139168 290898 139210 291134
rect 139446 290898 139488 291134
rect 139168 290866 139488 290898
rect 169888 291454 170208 291486
rect 169888 291218 169930 291454
rect 170166 291218 170208 291454
rect 169888 291134 170208 291218
rect 169888 290898 169930 291134
rect 170166 290898 170208 291134
rect 169888 290866 170208 290898
rect 200608 291454 200928 291486
rect 200608 291218 200650 291454
rect 200886 291218 200928 291454
rect 200608 291134 200928 291218
rect 200608 290898 200650 291134
rect 200886 290898 200928 291134
rect 200608 290866 200928 290898
rect 231328 291454 231648 291486
rect 231328 291218 231370 291454
rect 231606 291218 231648 291454
rect 231328 291134 231648 291218
rect 231328 290898 231370 291134
rect 231606 290898 231648 291134
rect 231328 290866 231648 290898
rect 262048 291454 262368 291486
rect 262048 291218 262090 291454
rect 262326 291218 262368 291454
rect 262048 291134 262368 291218
rect 262048 290898 262090 291134
rect 262326 290898 262368 291134
rect 262048 290866 262368 290898
rect 292768 291454 293088 291486
rect 292768 291218 292810 291454
rect 293046 291218 293088 291454
rect 292768 291134 293088 291218
rect 292768 290898 292810 291134
rect 293046 290898 293088 291134
rect 292768 290866 293088 290898
rect 323488 291454 323808 291486
rect 323488 291218 323530 291454
rect 323766 291218 323808 291454
rect 323488 291134 323808 291218
rect 323488 290898 323530 291134
rect 323766 290898 323808 291134
rect 323488 290866 323808 290898
rect 354208 291454 354528 291486
rect 354208 291218 354250 291454
rect 354486 291218 354528 291454
rect 354208 291134 354528 291218
rect 354208 290898 354250 291134
rect 354486 290898 354528 291134
rect 354208 290866 354528 290898
rect 384928 291454 385248 291486
rect 384928 291218 384970 291454
rect 385206 291218 385248 291454
rect 384928 291134 385248 291218
rect 384928 290898 384970 291134
rect 385206 290898 385248 291134
rect 384928 290866 385248 290898
rect 415648 291454 415968 291486
rect 415648 291218 415690 291454
rect 415926 291218 415968 291454
rect 415648 291134 415968 291218
rect 415648 290898 415690 291134
rect 415926 290898 415968 291134
rect 415648 290866 415968 290898
rect 446368 291454 446688 291486
rect 446368 291218 446410 291454
rect 446646 291218 446688 291454
rect 446368 291134 446688 291218
rect 446368 290898 446410 291134
rect 446646 290898 446688 291134
rect 446368 290866 446688 290898
rect 477088 291454 477408 291486
rect 477088 291218 477130 291454
rect 477366 291218 477408 291454
rect 477088 291134 477408 291218
rect 477088 290898 477130 291134
rect 477366 290898 477408 291134
rect 477088 290866 477408 290898
rect 507808 291454 508128 291486
rect 507808 291218 507850 291454
rect 508086 291218 508128 291454
rect 507808 291134 508128 291218
rect 507808 290898 507850 291134
rect 508086 290898 508128 291134
rect 507808 290866 508128 290898
rect 538528 291454 538848 291486
rect 538528 291218 538570 291454
rect 538806 291218 538848 291454
rect 538528 291134 538848 291218
rect 538528 290898 538570 291134
rect 538806 290898 538848 291134
rect 538528 290866 538848 290898
rect 62368 273454 62688 273486
rect 62368 273218 62410 273454
rect 62646 273218 62688 273454
rect 62368 273134 62688 273218
rect 62368 272898 62410 273134
rect 62646 272898 62688 273134
rect 62368 272866 62688 272898
rect 93088 273454 93408 273486
rect 93088 273218 93130 273454
rect 93366 273218 93408 273454
rect 93088 273134 93408 273218
rect 93088 272898 93130 273134
rect 93366 272898 93408 273134
rect 93088 272866 93408 272898
rect 123808 273454 124128 273486
rect 123808 273218 123850 273454
rect 124086 273218 124128 273454
rect 123808 273134 124128 273218
rect 123808 272898 123850 273134
rect 124086 272898 124128 273134
rect 123808 272866 124128 272898
rect 154528 273454 154848 273486
rect 154528 273218 154570 273454
rect 154806 273218 154848 273454
rect 154528 273134 154848 273218
rect 154528 272898 154570 273134
rect 154806 272898 154848 273134
rect 154528 272866 154848 272898
rect 185248 273454 185568 273486
rect 185248 273218 185290 273454
rect 185526 273218 185568 273454
rect 185248 273134 185568 273218
rect 185248 272898 185290 273134
rect 185526 272898 185568 273134
rect 185248 272866 185568 272898
rect 215968 273454 216288 273486
rect 215968 273218 216010 273454
rect 216246 273218 216288 273454
rect 215968 273134 216288 273218
rect 215968 272898 216010 273134
rect 216246 272898 216288 273134
rect 215968 272866 216288 272898
rect 246688 273454 247008 273486
rect 246688 273218 246730 273454
rect 246966 273218 247008 273454
rect 246688 273134 247008 273218
rect 246688 272898 246730 273134
rect 246966 272898 247008 273134
rect 246688 272866 247008 272898
rect 277408 273454 277728 273486
rect 277408 273218 277450 273454
rect 277686 273218 277728 273454
rect 277408 273134 277728 273218
rect 277408 272898 277450 273134
rect 277686 272898 277728 273134
rect 277408 272866 277728 272898
rect 308128 273454 308448 273486
rect 308128 273218 308170 273454
rect 308406 273218 308448 273454
rect 308128 273134 308448 273218
rect 308128 272898 308170 273134
rect 308406 272898 308448 273134
rect 308128 272866 308448 272898
rect 338848 273454 339168 273486
rect 338848 273218 338890 273454
rect 339126 273218 339168 273454
rect 338848 273134 339168 273218
rect 338848 272898 338890 273134
rect 339126 272898 339168 273134
rect 338848 272866 339168 272898
rect 369568 273454 369888 273486
rect 369568 273218 369610 273454
rect 369846 273218 369888 273454
rect 369568 273134 369888 273218
rect 369568 272898 369610 273134
rect 369846 272898 369888 273134
rect 369568 272866 369888 272898
rect 400288 273454 400608 273486
rect 400288 273218 400330 273454
rect 400566 273218 400608 273454
rect 400288 273134 400608 273218
rect 400288 272898 400330 273134
rect 400566 272898 400608 273134
rect 400288 272866 400608 272898
rect 431008 273454 431328 273486
rect 431008 273218 431050 273454
rect 431286 273218 431328 273454
rect 431008 273134 431328 273218
rect 431008 272898 431050 273134
rect 431286 272898 431328 273134
rect 431008 272866 431328 272898
rect 461728 273454 462048 273486
rect 461728 273218 461770 273454
rect 462006 273218 462048 273454
rect 461728 273134 462048 273218
rect 461728 272898 461770 273134
rect 462006 272898 462048 273134
rect 461728 272866 462048 272898
rect 492448 273454 492768 273486
rect 492448 273218 492490 273454
rect 492726 273218 492768 273454
rect 492448 273134 492768 273218
rect 492448 272898 492490 273134
rect 492726 272898 492768 273134
rect 492448 272866 492768 272898
rect 523168 273454 523488 273486
rect 523168 273218 523210 273454
rect 523446 273218 523488 273454
rect 523168 273134 523488 273218
rect 523168 272898 523210 273134
rect 523446 272898 523488 273134
rect 523168 272866 523488 272898
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 47008 255454 47328 255486
rect 47008 255218 47050 255454
rect 47286 255218 47328 255454
rect 47008 255134 47328 255218
rect 47008 254898 47050 255134
rect 47286 254898 47328 255134
rect 47008 254866 47328 254898
rect 77728 255454 78048 255486
rect 77728 255218 77770 255454
rect 78006 255218 78048 255454
rect 77728 255134 78048 255218
rect 77728 254898 77770 255134
rect 78006 254898 78048 255134
rect 77728 254866 78048 254898
rect 108448 255454 108768 255486
rect 108448 255218 108490 255454
rect 108726 255218 108768 255454
rect 108448 255134 108768 255218
rect 108448 254898 108490 255134
rect 108726 254898 108768 255134
rect 108448 254866 108768 254898
rect 139168 255454 139488 255486
rect 139168 255218 139210 255454
rect 139446 255218 139488 255454
rect 139168 255134 139488 255218
rect 139168 254898 139210 255134
rect 139446 254898 139488 255134
rect 139168 254866 139488 254898
rect 169888 255454 170208 255486
rect 169888 255218 169930 255454
rect 170166 255218 170208 255454
rect 169888 255134 170208 255218
rect 169888 254898 169930 255134
rect 170166 254898 170208 255134
rect 169888 254866 170208 254898
rect 200608 255454 200928 255486
rect 200608 255218 200650 255454
rect 200886 255218 200928 255454
rect 200608 255134 200928 255218
rect 200608 254898 200650 255134
rect 200886 254898 200928 255134
rect 200608 254866 200928 254898
rect 231328 255454 231648 255486
rect 231328 255218 231370 255454
rect 231606 255218 231648 255454
rect 231328 255134 231648 255218
rect 231328 254898 231370 255134
rect 231606 254898 231648 255134
rect 231328 254866 231648 254898
rect 262048 255454 262368 255486
rect 262048 255218 262090 255454
rect 262326 255218 262368 255454
rect 262048 255134 262368 255218
rect 262048 254898 262090 255134
rect 262326 254898 262368 255134
rect 262048 254866 262368 254898
rect 292768 255454 293088 255486
rect 292768 255218 292810 255454
rect 293046 255218 293088 255454
rect 292768 255134 293088 255218
rect 292768 254898 292810 255134
rect 293046 254898 293088 255134
rect 292768 254866 293088 254898
rect 323488 255454 323808 255486
rect 323488 255218 323530 255454
rect 323766 255218 323808 255454
rect 323488 255134 323808 255218
rect 323488 254898 323530 255134
rect 323766 254898 323808 255134
rect 323488 254866 323808 254898
rect 354208 255454 354528 255486
rect 354208 255218 354250 255454
rect 354486 255218 354528 255454
rect 354208 255134 354528 255218
rect 354208 254898 354250 255134
rect 354486 254898 354528 255134
rect 354208 254866 354528 254898
rect 384928 255454 385248 255486
rect 384928 255218 384970 255454
rect 385206 255218 385248 255454
rect 384928 255134 385248 255218
rect 384928 254898 384970 255134
rect 385206 254898 385248 255134
rect 384928 254866 385248 254898
rect 415648 255454 415968 255486
rect 415648 255218 415690 255454
rect 415926 255218 415968 255454
rect 415648 255134 415968 255218
rect 415648 254898 415690 255134
rect 415926 254898 415968 255134
rect 415648 254866 415968 254898
rect 446368 255454 446688 255486
rect 446368 255218 446410 255454
rect 446646 255218 446688 255454
rect 446368 255134 446688 255218
rect 446368 254898 446410 255134
rect 446646 254898 446688 255134
rect 446368 254866 446688 254898
rect 477088 255454 477408 255486
rect 477088 255218 477130 255454
rect 477366 255218 477408 255454
rect 477088 255134 477408 255218
rect 477088 254898 477130 255134
rect 477366 254898 477408 255134
rect 477088 254866 477408 254898
rect 507808 255454 508128 255486
rect 507808 255218 507850 255454
rect 508086 255218 508128 255454
rect 507808 255134 508128 255218
rect 507808 254898 507850 255134
rect 508086 254898 508128 255134
rect 507808 254866 508128 254898
rect 538528 255454 538848 255486
rect 538528 255218 538570 255454
rect 538806 255218 538848 255454
rect 538528 255134 538848 255218
rect 538528 254898 538570 255134
rect 538806 254898 538848 255134
rect 538528 254866 538848 254898
rect 62368 237454 62688 237486
rect 62368 237218 62410 237454
rect 62646 237218 62688 237454
rect 62368 237134 62688 237218
rect 62368 236898 62410 237134
rect 62646 236898 62688 237134
rect 62368 236866 62688 236898
rect 93088 237454 93408 237486
rect 93088 237218 93130 237454
rect 93366 237218 93408 237454
rect 93088 237134 93408 237218
rect 93088 236898 93130 237134
rect 93366 236898 93408 237134
rect 93088 236866 93408 236898
rect 123808 237454 124128 237486
rect 123808 237218 123850 237454
rect 124086 237218 124128 237454
rect 123808 237134 124128 237218
rect 123808 236898 123850 237134
rect 124086 236898 124128 237134
rect 123808 236866 124128 236898
rect 154528 237454 154848 237486
rect 154528 237218 154570 237454
rect 154806 237218 154848 237454
rect 154528 237134 154848 237218
rect 154528 236898 154570 237134
rect 154806 236898 154848 237134
rect 154528 236866 154848 236898
rect 185248 237454 185568 237486
rect 185248 237218 185290 237454
rect 185526 237218 185568 237454
rect 185248 237134 185568 237218
rect 185248 236898 185290 237134
rect 185526 236898 185568 237134
rect 185248 236866 185568 236898
rect 215968 237454 216288 237486
rect 215968 237218 216010 237454
rect 216246 237218 216288 237454
rect 215968 237134 216288 237218
rect 215968 236898 216010 237134
rect 216246 236898 216288 237134
rect 215968 236866 216288 236898
rect 246688 237454 247008 237486
rect 246688 237218 246730 237454
rect 246966 237218 247008 237454
rect 246688 237134 247008 237218
rect 246688 236898 246730 237134
rect 246966 236898 247008 237134
rect 246688 236866 247008 236898
rect 277408 237454 277728 237486
rect 277408 237218 277450 237454
rect 277686 237218 277728 237454
rect 277408 237134 277728 237218
rect 277408 236898 277450 237134
rect 277686 236898 277728 237134
rect 277408 236866 277728 236898
rect 308128 237454 308448 237486
rect 308128 237218 308170 237454
rect 308406 237218 308448 237454
rect 308128 237134 308448 237218
rect 308128 236898 308170 237134
rect 308406 236898 308448 237134
rect 308128 236866 308448 236898
rect 338848 237454 339168 237486
rect 338848 237218 338890 237454
rect 339126 237218 339168 237454
rect 338848 237134 339168 237218
rect 338848 236898 338890 237134
rect 339126 236898 339168 237134
rect 338848 236866 339168 236898
rect 369568 237454 369888 237486
rect 369568 237218 369610 237454
rect 369846 237218 369888 237454
rect 369568 237134 369888 237218
rect 369568 236898 369610 237134
rect 369846 236898 369888 237134
rect 369568 236866 369888 236898
rect 400288 237454 400608 237486
rect 400288 237218 400330 237454
rect 400566 237218 400608 237454
rect 400288 237134 400608 237218
rect 400288 236898 400330 237134
rect 400566 236898 400608 237134
rect 400288 236866 400608 236898
rect 431008 237454 431328 237486
rect 431008 237218 431050 237454
rect 431286 237218 431328 237454
rect 431008 237134 431328 237218
rect 431008 236898 431050 237134
rect 431286 236898 431328 237134
rect 431008 236866 431328 236898
rect 461728 237454 462048 237486
rect 461728 237218 461770 237454
rect 462006 237218 462048 237454
rect 461728 237134 462048 237218
rect 461728 236898 461770 237134
rect 462006 236898 462048 237134
rect 461728 236866 462048 236898
rect 492448 237454 492768 237486
rect 492448 237218 492490 237454
rect 492726 237218 492768 237454
rect 492448 237134 492768 237218
rect 492448 236898 492490 237134
rect 492726 236898 492768 237134
rect 492448 236866 492768 236898
rect 523168 237454 523488 237486
rect 523168 237218 523210 237454
rect 523446 237218 523488 237454
rect 523168 237134 523488 237218
rect 523168 236898 523210 237134
rect 523446 236898 523488 237134
rect 523168 236866 523488 236898
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 47008 219454 47328 219486
rect 47008 219218 47050 219454
rect 47286 219218 47328 219454
rect 47008 219134 47328 219218
rect 47008 218898 47050 219134
rect 47286 218898 47328 219134
rect 47008 218866 47328 218898
rect 77728 219454 78048 219486
rect 77728 219218 77770 219454
rect 78006 219218 78048 219454
rect 77728 219134 78048 219218
rect 77728 218898 77770 219134
rect 78006 218898 78048 219134
rect 77728 218866 78048 218898
rect 108448 219454 108768 219486
rect 108448 219218 108490 219454
rect 108726 219218 108768 219454
rect 108448 219134 108768 219218
rect 108448 218898 108490 219134
rect 108726 218898 108768 219134
rect 108448 218866 108768 218898
rect 139168 219454 139488 219486
rect 139168 219218 139210 219454
rect 139446 219218 139488 219454
rect 139168 219134 139488 219218
rect 139168 218898 139210 219134
rect 139446 218898 139488 219134
rect 139168 218866 139488 218898
rect 169888 219454 170208 219486
rect 169888 219218 169930 219454
rect 170166 219218 170208 219454
rect 169888 219134 170208 219218
rect 169888 218898 169930 219134
rect 170166 218898 170208 219134
rect 169888 218866 170208 218898
rect 200608 219454 200928 219486
rect 200608 219218 200650 219454
rect 200886 219218 200928 219454
rect 200608 219134 200928 219218
rect 200608 218898 200650 219134
rect 200886 218898 200928 219134
rect 200608 218866 200928 218898
rect 231328 219454 231648 219486
rect 231328 219218 231370 219454
rect 231606 219218 231648 219454
rect 231328 219134 231648 219218
rect 231328 218898 231370 219134
rect 231606 218898 231648 219134
rect 231328 218866 231648 218898
rect 262048 219454 262368 219486
rect 262048 219218 262090 219454
rect 262326 219218 262368 219454
rect 262048 219134 262368 219218
rect 262048 218898 262090 219134
rect 262326 218898 262368 219134
rect 262048 218866 262368 218898
rect 292768 219454 293088 219486
rect 292768 219218 292810 219454
rect 293046 219218 293088 219454
rect 292768 219134 293088 219218
rect 292768 218898 292810 219134
rect 293046 218898 293088 219134
rect 292768 218866 293088 218898
rect 323488 219454 323808 219486
rect 323488 219218 323530 219454
rect 323766 219218 323808 219454
rect 323488 219134 323808 219218
rect 323488 218898 323530 219134
rect 323766 218898 323808 219134
rect 323488 218866 323808 218898
rect 354208 219454 354528 219486
rect 354208 219218 354250 219454
rect 354486 219218 354528 219454
rect 354208 219134 354528 219218
rect 354208 218898 354250 219134
rect 354486 218898 354528 219134
rect 354208 218866 354528 218898
rect 384928 219454 385248 219486
rect 384928 219218 384970 219454
rect 385206 219218 385248 219454
rect 384928 219134 385248 219218
rect 384928 218898 384970 219134
rect 385206 218898 385248 219134
rect 384928 218866 385248 218898
rect 415648 219454 415968 219486
rect 415648 219218 415690 219454
rect 415926 219218 415968 219454
rect 415648 219134 415968 219218
rect 415648 218898 415690 219134
rect 415926 218898 415968 219134
rect 415648 218866 415968 218898
rect 446368 219454 446688 219486
rect 446368 219218 446410 219454
rect 446646 219218 446688 219454
rect 446368 219134 446688 219218
rect 446368 218898 446410 219134
rect 446646 218898 446688 219134
rect 446368 218866 446688 218898
rect 477088 219454 477408 219486
rect 477088 219218 477130 219454
rect 477366 219218 477408 219454
rect 477088 219134 477408 219218
rect 477088 218898 477130 219134
rect 477366 218898 477408 219134
rect 477088 218866 477408 218898
rect 507808 219454 508128 219486
rect 507808 219218 507850 219454
rect 508086 219218 508128 219454
rect 507808 219134 508128 219218
rect 507808 218898 507850 219134
rect 508086 218898 508128 219134
rect 507808 218866 508128 218898
rect 538528 219454 538848 219486
rect 538528 219218 538570 219454
rect 538806 219218 538848 219454
rect 538528 219134 538848 219218
rect 538528 218898 538570 219134
rect 538806 218898 538848 219134
rect 538528 218866 538848 218898
rect 62368 201454 62688 201486
rect 62368 201218 62410 201454
rect 62646 201218 62688 201454
rect 62368 201134 62688 201218
rect 62368 200898 62410 201134
rect 62646 200898 62688 201134
rect 62368 200866 62688 200898
rect 93088 201454 93408 201486
rect 93088 201218 93130 201454
rect 93366 201218 93408 201454
rect 93088 201134 93408 201218
rect 93088 200898 93130 201134
rect 93366 200898 93408 201134
rect 93088 200866 93408 200898
rect 123808 201454 124128 201486
rect 123808 201218 123850 201454
rect 124086 201218 124128 201454
rect 123808 201134 124128 201218
rect 123808 200898 123850 201134
rect 124086 200898 124128 201134
rect 123808 200866 124128 200898
rect 154528 201454 154848 201486
rect 154528 201218 154570 201454
rect 154806 201218 154848 201454
rect 154528 201134 154848 201218
rect 154528 200898 154570 201134
rect 154806 200898 154848 201134
rect 154528 200866 154848 200898
rect 185248 201454 185568 201486
rect 185248 201218 185290 201454
rect 185526 201218 185568 201454
rect 185248 201134 185568 201218
rect 185248 200898 185290 201134
rect 185526 200898 185568 201134
rect 185248 200866 185568 200898
rect 215968 201454 216288 201486
rect 215968 201218 216010 201454
rect 216246 201218 216288 201454
rect 215968 201134 216288 201218
rect 215968 200898 216010 201134
rect 216246 200898 216288 201134
rect 215968 200866 216288 200898
rect 246688 201454 247008 201486
rect 246688 201218 246730 201454
rect 246966 201218 247008 201454
rect 246688 201134 247008 201218
rect 246688 200898 246730 201134
rect 246966 200898 247008 201134
rect 246688 200866 247008 200898
rect 277408 201454 277728 201486
rect 277408 201218 277450 201454
rect 277686 201218 277728 201454
rect 277408 201134 277728 201218
rect 277408 200898 277450 201134
rect 277686 200898 277728 201134
rect 277408 200866 277728 200898
rect 308128 201454 308448 201486
rect 308128 201218 308170 201454
rect 308406 201218 308448 201454
rect 308128 201134 308448 201218
rect 308128 200898 308170 201134
rect 308406 200898 308448 201134
rect 308128 200866 308448 200898
rect 338848 201454 339168 201486
rect 338848 201218 338890 201454
rect 339126 201218 339168 201454
rect 338848 201134 339168 201218
rect 338848 200898 338890 201134
rect 339126 200898 339168 201134
rect 338848 200866 339168 200898
rect 369568 201454 369888 201486
rect 369568 201218 369610 201454
rect 369846 201218 369888 201454
rect 369568 201134 369888 201218
rect 369568 200898 369610 201134
rect 369846 200898 369888 201134
rect 369568 200866 369888 200898
rect 400288 201454 400608 201486
rect 400288 201218 400330 201454
rect 400566 201218 400608 201454
rect 400288 201134 400608 201218
rect 400288 200898 400330 201134
rect 400566 200898 400608 201134
rect 400288 200866 400608 200898
rect 431008 201454 431328 201486
rect 431008 201218 431050 201454
rect 431286 201218 431328 201454
rect 431008 201134 431328 201218
rect 431008 200898 431050 201134
rect 431286 200898 431328 201134
rect 431008 200866 431328 200898
rect 461728 201454 462048 201486
rect 461728 201218 461770 201454
rect 462006 201218 462048 201454
rect 461728 201134 462048 201218
rect 461728 200898 461770 201134
rect 462006 200898 462048 201134
rect 461728 200866 462048 200898
rect 492448 201454 492768 201486
rect 492448 201218 492490 201454
rect 492726 201218 492768 201454
rect 492448 201134 492768 201218
rect 492448 200898 492490 201134
rect 492726 200898 492768 201134
rect 492448 200866 492768 200898
rect 523168 201454 523488 201486
rect 523168 201218 523210 201454
rect 523446 201218 523488 201454
rect 523168 201134 523488 201218
rect 523168 200898 523210 201134
rect 523446 200898 523488 201134
rect 523168 200866 523488 200898
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 47008 183454 47328 183486
rect 47008 183218 47050 183454
rect 47286 183218 47328 183454
rect 47008 183134 47328 183218
rect 47008 182898 47050 183134
rect 47286 182898 47328 183134
rect 47008 182866 47328 182898
rect 77728 183454 78048 183486
rect 77728 183218 77770 183454
rect 78006 183218 78048 183454
rect 77728 183134 78048 183218
rect 77728 182898 77770 183134
rect 78006 182898 78048 183134
rect 77728 182866 78048 182898
rect 108448 183454 108768 183486
rect 108448 183218 108490 183454
rect 108726 183218 108768 183454
rect 108448 183134 108768 183218
rect 108448 182898 108490 183134
rect 108726 182898 108768 183134
rect 108448 182866 108768 182898
rect 139168 183454 139488 183486
rect 139168 183218 139210 183454
rect 139446 183218 139488 183454
rect 139168 183134 139488 183218
rect 139168 182898 139210 183134
rect 139446 182898 139488 183134
rect 139168 182866 139488 182898
rect 169888 183454 170208 183486
rect 169888 183218 169930 183454
rect 170166 183218 170208 183454
rect 169888 183134 170208 183218
rect 169888 182898 169930 183134
rect 170166 182898 170208 183134
rect 169888 182866 170208 182898
rect 200608 183454 200928 183486
rect 200608 183218 200650 183454
rect 200886 183218 200928 183454
rect 200608 183134 200928 183218
rect 200608 182898 200650 183134
rect 200886 182898 200928 183134
rect 200608 182866 200928 182898
rect 231328 183454 231648 183486
rect 231328 183218 231370 183454
rect 231606 183218 231648 183454
rect 231328 183134 231648 183218
rect 231328 182898 231370 183134
rect 231606 182898 231648 183134
rect 231328 182866 231648 182898
rect 262048 183454 262368 183486
rect 262048 183218 262090 183454
rect 262326 183218 262368 183454
rect 262048 183134 262368 183218
rect 262048 182898 262090 183134
rect 262326 182898 262368 183134
rect 262048 182866 262368 182898
rect 292768 183454 293088 183486
rect 292768 183218 292810 183454
rect 293046 183218 293088 183454
rect 292768 183134 293088 183218
rect 292768 182898 292810 183134
rect 293046 182898 293088 183134
rect 292768 182866 293088 182898
rect 323488 183454 323808 183486
rect 323488 183218 323530 183454
rect 323766 183218 323808 183454
rect 323488 183134 323808 183218
rect 323488 182898 323530 183134
rect 323766 182898 323808 183134
rect 323488 182866 323808 182898
rect 354208 183454 354528 183486
rect 354208 183218 354250 183454
rect 354486 183218 354528 183454
rect 354208 183134 354528 183218
rect 354208 182898 354250 183134
rect 354486 182898 354528 183134
rect 354208 182866 354528 182898
rect 384928 183454 385248 183486
rect 384928 183218 384970 183454
rect 385206 183218 385248 183454
rect 384928 183134 385248 183218
rect 384928 182898 384970 183134
rect 385206 182898 385248 183134
rect 384928 182866 385248 182898
rect 415648 183454 415968 183486
rect 415648 183218 415690 183454
rect 415926 183218 415968 183454
rect 415648 183134 415968 183218
rect 415648 182898 415690 183134
rect 415926 182898 415968 183134
rect 415648 182866 415968 182898
rect 446368 183454 446688 183486
rect 446368 183218 446410 183454
rect 446646 183218 446688 183454
rect 446368 183134 446688 183218
rect 446368 182898 446410 183134
rect 446646 182898 446688 183134
rect 446368 182866 446688 182898
rect 477088 183454 477408 183486
rect 477088 183218 477130 183454
rect 477366 183218 477408 183454
rect 477088 183134 477408 183218
rect 477088 182898 477130 183134
rect 477366 182898 477408 183134
rect 477088 182866 477408 182898
rect 507808 183454 508128 183486
rect 507808 183218 507850 183454
rect 508086 183218 508128 183454
rect 507808 183134 508128 183218
rect 507808 182898 507850 183134
rect 508086 182898 508128 183134
rect 507808 182866 508128 182898
rect 538528 183454 538848 183486
rect 538528 183218 538570 183454
rect 538806 183218 538848 183454
rect 538528 183134 538848 183218
rect 538528 182898 538570 183134
rect 538806 182898 538848 183134
rect 538528 182866 538848 182898
rect 62368 165454 62688 165486
rect 62368 165218 62410 165454
rect 62646 165218 62688 165454
rect 62368 165134 62688 165218
rect 62368 164898 62410 165134
rect 62646 164898 62688 165134
rect 62368 164866 62688 164898
rect 93088 165454 93408 165486
rect 93088 165218 93130 165454
rect 93366 165218 93408 165454
rect 93088 165134 93408 165218
rect 93088 164898 93130 165134
rect 93366 164898 93408 165134
rect 93088 164866 93408 164898
rect 123808 165454 124128 165486
rect 123808 165218 123850 165454
rect 124086 165218 124128 165454
rect 123808 165134 124128 165218
rect 123808 164898 123850 165134
rect 124086 164898 124128 165134
rect 123808 164866 124128 164898
rect 154528 165454 154848 165486
rect 154528 165218 154570 165454
rect 154806 165218 154848 165454
rect 154528 165134 154848 165218
rect 154528 164898 154570 165134
rect 154806 164898 154848 165134
rect 154528 164866 154848 164898
rect 185248 165454 185568 165486
rect 185248 165218 185290 165454
rect 185526 165218 185568 165454
rect 185248 165134 185568 165218
rect 185248 164898 185290 165134
rect 185526 164898 185568 165134
rect 185248 164866 185568 164898
rect 215968 165454 216288 165486
rect 215968 165218 216010 165454
rect 216246 165218 216288 165454
rect 215968 165134 216288 165218
rect 215968 164898 216010 165134
rect 216246 164898 216288 165134
rect 215968 164866 216288 164898
rect 246688 165454 247008 165486
rect 246688 165218 246730 165454
rect 246966 165218 247008 165454
rect 246688 165134 247008 165218
rect 246688 164898 246730 165134
rect 246966 164898 247008 165134
rect 246688 164866 247008 164898
rect 277408 165454 277728 165486
rect 277408 165218 277450 165454
rect 277686 165218 277728 165454
rect 277408 165134 277728 165218
rect 277408 164898 277450 165134
rect 277686 164898 277728 165134
rect 277408 164866 277728 164898
rect 308128 165454 308448 165486
rect 308128 165218 308170 165454
rect 308406 165218 308448 165454
rect 308128 165134 308448 165218
rect 308128 164898 308170 165134
rect 308406 164898 308448 165134
rect 308128 164866 308448 164898
rect 338848 165454 339168 165486
rect 338848 165218 338890 165454
rect 339126 165218 339168 165454
rect 338848 165134 339168 165218
rect 338848 164898 338890 165134
rect 339126 164898 339168 165134
rect 338848 164866 339168 164898
rect 369568 165454 369888 165486
rect 369568 165218 369610 165454
rect 369846 165218 369888 165454
rect 369568 165134 369888 165218
rect 369568 164898 369610 165134
rect 369846 164898 369888 165134
rect 369568 164866 369888 164898
rect 400288 165454 400608 165486
rect 400288 165218 400330 165454
rect 400566 165218 400608 165454
rect 400288 165134 400608 165218
rect 400288 164898 400330 165134
rect 400566 164898 400608 165134
rect 400288 164866 400608 164898
rect 431008 165454 431328 165486
rect 431008 165218 431050 165454
rect 431286 165218 431328 165454
rect 431008 165134 431328 165218
rect 431008 164898 431050 165134
rect 431286 164898 431328 165134
rect 431008 164866 431328 164898
rect 461728 165454 462048 165486
rect 461728 165218 461770 165454
rect 462006 165218 462048 165454
rect 461728 165134 462048 165218
rect 461728 164898 461770 165134
rect 462006 164898 462048 165134
rect 461728 164866 462048 164898
rect 492448 165454 492768 165486
rect 492448 165218 492490 165454
rect 492726 165218 492768 165454
rect 492448 165134 492768 165218
rect 492448 164898 492490 165134
rect 492726 164898 492768 165134
rect 492448 164866 492768 164898
rect 523168 165454 523488 165486
rect 523168 165218 523210 165454
rect 523446 165218 523488 165454
rect 523168 165134 523488 165218
rect 523168 164898 523210 165134
rect 523446 164898 523488 165134
rect 523168 164866 523488 164898
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 47008 147454 47328 147486
rect 47008 147218 47050 147454
rect 47286 147218 47328 147454
rect 47008 147134 47328 147218
rect 47008 146898 47050 147134
rect 47286 146898 47328 147134
rect 47008 146866 47328 146898
rect 77728 147454 78048 147486
rect 77728 147218 77770 147454
rect 78006 147218 78048 147454
rect 77728 147134 78048 147218
rect 77728 146898 77770 147134
rect 78006 146898 78048 147134
rect 77728 146866 78048 146898
rect 108448 147454 108768 147486
rect 108448 147218 108490 147454
rect 108726 147218 108768 147454
rect 108448 147134 108768 147218
rect 108448 146898 108490 147134
rect 108726 146898 108768 147134
rect 108448 146866 108768 146898
rect 139168 147454 139488 147486
rect 139168 147218 139210 147454
rect 139446 147218 139488 147454
rect 139168 147134 139488 147218
rect 139168 146898 139210 147134
rect 139446 146898 139488 147134
rect 139168 146866 139488 146898
rect 169888 147454 170208 147486
rect 169888 147218 169930 147454
rect 170166 147218 170208 147454
rect 169888 147134 170208 147218
rect 169888 146898 169930 147134
rect 170166 146898 170208 147134
rect 169888 146866 170208 146898
rect 200608 147454 200928 147486
rect 200608 147218 200650 147454
rect 200886 147218 200928 147454
rect 200608 147134 200928 147218
rect 200608 146898 200650 147134
rect 200886 146898 200928 147134
rect 200608 146866 200928 146898
rect 231328 147454 231648 147486
rect 231328 147218 231370 147454
rect 231606 147218 231648 147454
rect 231328 147134 231648 147218
rect 231328 146898 231370 147134
rect 231606 146898 231648 147134
rect 231328 146866 231648 146898
rect 262048 147454 262368 147486
rect 262048 147218 262090 147454
rect 262326 147218 262368 147454
rect 262048 147134 262368 147218
rect 262048 146898 262090 147134
rect 262326 146898 262368 147134
rect 262048 146866 262368 146898
rect 292768 147454 293088 147486
rect 292768 147218 292810 147454
rect 293046 147218 293088 147454
rect 292768 147134 293088 147218
rect 292768 146898 292810 147134
rect 293046 146898 293088 147134
rect 292768 146866 293088 146898
rect 323488 147454 323808 147486
rect 323488 147218 323530 147454
rect 323766 147218 323808 147454
rect 323488 147134 323808 147218
rect 323488 146898 323530 147134
rect 323766 146898 323808 147134
rect 323488 146866 323808 146898
rect 354208 147454 354528 147486
rect 354208 147218 354250 147454
rect 354486 147218 354528 147454
rect 354208 147134 354528 147218
rect 354208 146898 354250 147134
rect 354486 146898 354528 147134
rect 354208 146866 354528 146898
rect 384928 147454 385248 147486
rect 384928 147218 384970 147454
rect 385206 147218 385248 147454
rect 384928 147134 385248 147218
rect 384928 146898 384970 147134
rect 385206 146898 385248 147134
rect 384928 146866 385248 146898
rect 415648 147454 415968 147486
rect 415648 147218 415690 147454
rect 415926 147218 415968 147454
rect 415648 147134 415968 147218
rect 415648 146898 415690 147134
rect 415926 146898 415968 147134
rect 415648 146866 415968 146898
rect 446368 147454 446688 147486
rect 446368 147218 446410 147454
rect 446646 147218 446688 147454
rect 446368 147134 446688 147218
rect 446368 146898 446410 147134
rect 446646 146898 446688 147134
rect 446368 146866 446688 146898
rect 477088 147454 477408 147486
rect 477088 147218 477130 147454
rect 477366 147218 477408 147454
rect 477088 147134 477408 147218
rect 477088 146898 477130 147134
rect 477366 146898 477408 147134
rect 477088 146866 477408 146898
rect 507808 147454 508128 147486
rect 507808 147218 507850 147454
rect 508086 147218 508128 147454
rect 507808 147134 508128 147218
rect 507808 146898 507850 147134
rect 508086 146898 508128 147134
rect 507808 146866 508128 146898
rect 538528 147454 538848 147486
rect 538528 147218 538570 147454
rect 538806 147218 538848 147454
rect 538528 147134 538848 147218
rect 538528 146898 538570 147134
rect 538806 146898 538848 147134
rect 538528 146866 538848 146898
rect 62368 129454 62688 129486
rect 62368 129218 62410 129454
rect 62646 129218 62688 129454
rect 62368 129134 62688 129218
rect 62368 128898 62410 129134
rect 62646 128898 62688 129134
rect 62368 128866 62688 128898
rect 93088 129454 93408 129486
rect 93088 129218 93130 129454
rect 93366 129218 93408 129454
rect 93088 129134 93408 129218
rect 93088 128898 93130 129134
rect 93366 128898 93408 129134
rect 93088 128866 93408 128898
rect 123808 129454 124128 129486
rect 123808 129218 123850 129454
rect 124086 129218 124128 129454
rect 123808 129134 124128 129218
rect 123808 128898 123850 129134
rect 124086 128898 124128 129134
rect 123808 128866 124128 128898
rect 154528 129454 154848 129486
rect 154528 129218 154570 129454
rect 154806 129218 154848 129454
rect 154528 129134 154848 129218
rect 154528 128898 154570 129134
rect 154806 128898 154848 129134
rect 154528 128866 154848 128898
rect 185248 129454 185568 129486
rect 185248 129218 185290 129454
rect 185526 129218 185568 129454
rect 185248 129134 185568 129218
rect 185248 128898 185290 129134
rect 185526 128898 185568 129134
rect 185248 128866 185568 128898
rect 215968 129454 216288 129486
rect 215968 129218 216010 129454
rect 216246 129218 216288 129454
rect 215968 129134 216288 129218
rect 215968 128898 216010 129134
rect 216246 128898 216288 129134
rect 215968 128866 216288 128898
rect 246688 129454 247008 129486
rect 246688 129218 246730 129454
rect 246966 129218 247008 129454
rect 246688 129134 247008 129218
rect 246688 128898 246730 129134
rect 246966 128898 247008 129134
rect 246688 128866 247008 128898
rect 277408 129454 277728 129486
rect 277408 129218 277450 129454
rect 277686 129218 277728 129454
rect 277408 129134 277728 129218
rect 277408 128898 277450 129134
rect 277686 128898 277728 129134
rect 277408 128866 277728 128898
rect 308128 129454 308448 129486
rect 308128 129218 308170 129454
rect 308406 129218 308448 129454
rect 308128 129134 308448 129218
rect 308128 128898 308170 129134
rect 308406 128898 308448 129134
rect 308128 128866 308448 128898
rect 338848 129454 339168 129486
rect 338848 129218 338890 129454
rect 339126 129218 339168 129454
rect 338848 129134 339168 129218
rect 338848 128898 338890 129134
rect 339126 128898 339168 129134
rect 338848 128866 339168 128898
rect 369568 129454 369888 129486
rect 369568 129218 369610 129454
rect 369846 129218 369888 129454
rect 369568 129134 369888 129218
rect 369568 128898 369610 129134
rect 369846 128898 369888 129134
rect 369568 128866 369888 128898
rect 400288 129454 400608 129486
rect 400288 129218 400330 129454
rect 400566 129218 400608 129454
rect 400288 129134 400608 129218
rect 400288 128898 400330 129134
rect 400566 128898 400608 129134
rect 400288 128866 400608 128898
rect 431008 129454 431328 129486
rect 431008 129218 431050 129454
rect 431286 129218 431328 129454
rect 431008 129134 431328 129218
rect 431008 128898 431050 129134
rect 431286 128898 431328 129134
rect 431008 128866 431328 128898
rect 461728 129454 462048 129486
rect 461728 129218 461770 129454
rect 462006 129218 462048 129454
rect 461728 129134 462048 129218
rect 461728 128898 461770 129134
rect 462006 128898 462048 129134
rect 461728 128866 462048 128898
rect 492448 129454 492768 129486
rect 492448 129218 492490 129454
rect 492726 129218 492768 129454
rect 492448 129134 492768 129218
rect 492448 128898 492490 129134
rect 492726 128898 492768 129134
rect 492448 128866 492768 128898
rect 523168 129454 523488 129486
rect 523168 129218 523210 129454
rect 523446 129218 523488 129454
rect 523168 129134 523488 129218
rect 523168 128898 523210 129134
rect 523446 128898 523488 129134
rect 523168 128866 523488 128898
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 47008 111454 47328 111486
rect 47008 111218 47050 111454
rect 47286 111218 47328 111454
rect 47008 111134 47328 111218
rect 47008 110898 47050 111134
rect 47286 110898 47328 111134
rect 47008 110866 47328 110898
rect 77728 111454 78048 111486
rect 77728 111218 77770 111454
rect 78006 111218 78048 111454
rect 77728 111134 78048 111218
rect 77728 110898 77770 111134
rect 78006 110898 78048 111134
rect 77728 110866 78048 110898
rect 108448 111454 108768 111486
rect 108448 111218 108490 111454
rect 108726 111218 108768 111454
rect 108448 111134 108768 111218
rect 108448 110898 108490 111134
rect 108726 110898 108768 111134
rect 108448 110866 108768 110898
rect 139168 111454 139488 111486
rect 139168 111218 139210 111454
rect 139446 111218 139488 111454
rect 139168 111134 139488 111218
rect 139168 110898 139210 111134
rect 139446 110898 139488 111134
rect 139168 110866 139488 110898
rect 169888 111454 170208 111486
rect 169888 111218 169930 111454
rect 170166 111218 170208 111454
rect 169888 111134 170208 111218
rect 169888 110898 169930 111134
rect 170166 110898 170208 111134
rect 169888 110866 170208 110898
rect 200608 111454 200928 111486
rect 200608 111218 200650 111454
rect 200886 111218 200928 111454
rect 200608 111134 200928 111218
rect 200608 110898 200650 111134
rect 200886 110898 200928 111134
rect 200608 110866 200928 110898
rect 231328 111454 231648 111486
rect 231328 111218 231370 111454
rect 231606 111218 231648 111454
rect 231328 111134 231648 111218
rect 231328 110898 231370 111134
rect 231606 110898 231648 111134
rect 231328 110866 231648 110898
rect 262048 111454 262368 111486
rect 262048 111218 262090 111454
rect 262326 111218 262368 111454
rect 262048 111134 262368 111218
rect 262048 110898 262090 111134
rect 262326 110898 262368 111134
rect 262048 110866 262368 110898
rect 292768 111454 293088 111486
rect 292768 111218 292810 111454
rect 293046 111218 293088 111454
rect 292768 111134 293088 111218
rect 292768 110898 292810 111134
rect 293046 110898 293088 111134
rect 292768 110866 293088 110898
rect 323488 111454 323808 111486
rect 323488 111218 323530 111454
rect 323766 111218 323808 111454
rect 323488 111134 323808 111218
rect 323488 110898 323530 111134
rect 323766 110898 323808 111134
rect 323488 110866 323808 110898
rect 354208 111454 354528 111486
rect 354208 111218 354250 111454
rect 354486 111218 354528 111454
rect 354208 111134 354528 111218
rect 354208 110898 354250 111134
rect 354486 110898 354528 111134
rect 354208 110866 354528 110898
rect 384928 111454 385248 111486
rect 384928 111218 384970 111454
rect 385206 111218 385248 111454
rect 384928 111134 385248 111218
rect 384928 110898 384970 111134
rect 385206 110898 385248 111134
rect 384928 110866 385248 110898
rect 415648 111454 415968 111486
rect 415648 111218 415690 111454
rect 415926 111218 415968 111454
rect 415648 111134 415968 111218
rect 415648 110898 415690 111134
rect 415926 110898 415968 111134
rect 415648 110866 415968 110898
rect 446368 111454 446688 111486
rect 446368 111218 446410 111454
rect 446646 111218 446688 111454
rect 446368 111134 446688 111218
rect 446368 110898 446410 111134
rect 446646 110898 446688 111134
rect 446368 110866 446688 110898
rect 477088 111454 477408 111486
rect 477088 111218 477130 111454
rect 477366 111218 477408 111454
rect 477088 111134 477408 111218
rect 477088 110898 477130 111134
rect 477366 110898 477408 111134
rect 477088 110866 477408 110898
rect 507808 111454 508128 111486
rect 507808 111218 507850 111454
rect 508086 111218 508128 111454
rect 507808 111134 508128 111218
rect 507808 110898 507850 111134
rect 508086 110898 508128 111134
rect 507808 110866 508128 110898
rect 538528 111454 538848 111486
rect 538528 111218 538570 111454
rect 538806 111218 538848 111454
rect 538528 111134 538848 111218
rect 538528 110898 538570 111134
rect 538806 110898 538848 111134
rect 538528 110866 538848 110898
rect 62368 93454 62688 93486
rect 62368 93218 62410 93454
rect 62646 93218 62688 93454
rect 62368 93134 62688 93218
rect 62368 92898 62410 93134
rect 62646 92898 62688 93134
rect 62368 92866 62688 92898
rect 93088 93454 93408 93486
rect 93088 93218 93130 93454
rect 93366 93218 93408 93454
rect 93088 93134 93408 93218
rect 93088 92898 93130 93134
rect 93366 92898 93408 93134
rect 93088 92866 93408 92898
rect 123808 93454 124128 93486
rect 123808 93218 123850 93454
rect 124086 93218 124128 93454
rect 123808 93134 124128 93218
rect 123808 92898 123850 93134
rect 124086 92898 124128 93134
rect 123808 92866 124128 92898
rect 154528 93454 154848 93486
rect 154528 93218 154570 93454
rect 154806 93218 154848 93454
rect 154528 93134 154848 93218
rect 154528 92898 154570 93134
rect 154806 92898 154848 93134
rect 154528 92866 154848 92898
rect 185248 93454 185568 93486
rect 185248 93218 185290 93454
rect 185526 93218 185568 93454
rect 185248 93134 185568 93218
rect 185248 92898 185290 93134
rect 185526 92898 185568 93134
rect 185248 92866 185568 92898
rect 215968 93454 216288 93486
rect 215968 93218 216010 93454
rect 216246 93218 216288 93454
rect 215968 93134 216288 93218
rect 215968 92898 216010 93134
rect 216246 92898 216288 93134
rect 215968 92866 216288 92898
rect 246688 93454 247008 93486
rect 246688 93218 246730 93454
rect 246966 93218 247008 93454
rect 246688 93134 247008 93218
rect 246688 92898 246730 93134
rect 246966 92898 247008 93134
rect 246688 92866 247008 92898
rect 277408 93454 277728 93486
rect 277408 93218 277450 93454
rect 277686 93218 277728 93454
rect 277408 93134 277728 93218
rect 277408 92898 277450 93134
rect 277686 92898 277728 93134
rect 277408 92866 277728 92898
rect 308128 93454 308448 93486
rect 308128 93218 308170 93454
rect 308406 93218 308448 93454
rect 308128 93134 308448 93218
rect 308128 92898 308170 93134
rect 308406 92898 308448 93134
rect 308128 92866 308448 92898
rect 338848 93454 339168 93486
rect 338848 93218 338890 93454
rect 339126 93218 339168 93454
rect 338848 93134 339168 93218
rect 338848 92898 338890 93134
rect 339126 92898 339168 93134
rect 338848 92866 339168 92898
rect 369568 93454 369888 93486
rect 369568 93218 369610 93454
rect 369846 93218 369888 93454
rect 369568 93134 369888 93218
rect 369568 92898 369610 93134
rect 369846 92898 369888 93134
rect 369568 92866 369888 92898
rect 400288 93454 400608 93486
rect 400288 93218 400330 93454
rect 400566 93218 400608 93454
rect 400288 93134 400608 93218
rect 400288 92898 400330 93134
rect 400566 92898 400608 93134
rect 400288 92866 400608 92898
rect 431008 93454 431328 93486
rect 431008 93218 431050 93454
rect 431286 93218 431328 93454
rect 431008 93134 431328 93218
rect 431008 92898 431050 93134
rect 431286 92898 431328 93134
rect 431008 92866 431328 92898
rect 461728 93454 462048 93486
rect 461728 93218 461770 93454
rect 462006 93218 462048 93454
rect 461728 93134 462048 93218
rect 461728 92898 461770 93134
rect 462006 92898 462048 93134
rect 461728 92866 462048 92898
rect 492448 93454 492768 93486
rect 492448 93218 492490 93454
rect 492726 93218 492768 93454
rect 492448 93134 492768 93218
rect 492448 92898 492490 93134
rect 492726 92898 492768 93134
rect 492448 92866 492768 92898
rect 523168 93454 523488 93486
rect 523168 93218 523210 93454
rect 523446 93218 523488 93454
rect 523168 93134 523488 93218
rect 523168 92898 523210 93134
rect 523446 92898 523488 93134
rect 523168 92866 523488 92898
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 47008 75454 47328 75486
rect 47008 75218 47050 75454
rect 47286 75218 47328 75454
rect 47008 75134 47328 75218
rect 47008 74898 47050 75134
rect 47286 74898 47328 75134
rect 47008 74866 47328 74898
rect 77728 75454 78048 75486
rect 77728 75218 77770 75454
rect 78006 75218 78048 75454
rect 77728 75134 78048 75218
rect 77728 74898 77770 75134
rect 78006 74898 78048 75134
rect 77728 74866 78048 74898
rect 108448 75454 108768 75486
rect 108448 75218 108490 75454
rect 108726 75218 108768 75454
rect 108448 75134 108768 75218
rect 108448 74898 108490 75134
rect 108726 74898 108768 75134
rect 108448 74866 108768 74898
rect 139168 75454 139488 75486
rect 139168 75218 139210 75454
rect 139446 75218 139488 75454
rect 139168 75134 139488 75218
rect 139168 74898 139210 75134
rect 139446 74898 139488 75134
rect 139168 74866 139488 74898
rect 169888 75454 170208 75486
rect 169888 75218 169930 75454
rect 170166 75218 170208 75454
rect 169888 75134 170208 75218
rect 169888 74898 169930 75134
rect 170166 74898 170208 75134
rect 169888 74866 170208 74898
rect 200608 75454 200928 75486
rect 200608 75218 200650 75454
rect 200886 75218 200928 75454
rect 200608 75134 200928 75218
rect 200608 74898 200650 75134
rect 200886 74898 200928 75134
rect 200608 74866 200928 74898
rect 231328 75454 231648 75486
rect 231328 75218 231370 75454
rect 231606 75218 231648 75454
rect 231328 75134 231648 75218
rect 231328 74898 231370 75134
rect 231606 74898 231648 75134
rect 231328 74866 231648 74898
rect 262048 75454 262368 75486
rect 262048 75218 262090 75454
rect 262326 75218 262368 75454
rect 262048 75134 262368 75218
rect 262048 74898 262090 75134
rect 262326 74898 262368 75134
rect 262048 74866 262368 74898
rect 292768 75454 293088 75486
rect 292768 75218 292810 75454
rect 293046 75218 293088 75454
rect 292768 75134 293088 75218
rect 292768 74898 292810 75134
rect 293046 74898 293088 75134
rect 292768 74866 293088 74898
rect 323488 75454 323808 75486
rect 323488 75218 323530 75454
rect 323766 75218 323808 75454
rect 323488 75134 323808 75218
rect 323488 74898 323530 75134
rect 323766 74898 323808 75134
rect 323488 74866 323808 74898
rect 354208 75454 354528 75486
rect 354208 75218 354250 75454
rect 354486 75218 354528 75454
rect 354208 75134 354528 75218
rect 354208 74898 354250 75134
rect 354486 74898 354528 75134
rect 354208 74866 354528 74898
rect 384928 75454 385248 75486
rect 384928 75218 384970 75454
rect 385206 75218 385248 75454
rect 384928 75134 385248 75218
rect 384928 74898 384970 75134
rect 385206 74898 385248 75134
rect 384928 74866 385248 74898
rect 415648 75454 415968 75486
rect 415648 75218 415690 75454
rect 415926 75218 415968 75454
rect 415648 75134 415968 75218
rect 415648 74898 415690 75134
rect 415926 74898 415968 75134
rect 415648 74866 415968 74898
rect 446368 75454 446688 75486
rect 446368 75218 446410 75454
rect 446646 75218 446688 75454
rect 446368 75134 446688 75218
rect 446368 74898 446410 75134
rect 446646 74898 446688 75134
rect 446368 74866 446688 74898
rect 477088 75454 477408 75486
rect 477088 75218 477130 75454
rect 477366 75218 477408 75454
rect 477088 75134 477408 75218
rect 477088 74898 477130 75134
rect 477366 74898 477408 75134
rect 477088 74866 477408 74898
rect 507808 75454 508128 75486
rect 507808 75218 507850 75454
rect 508086 75218 508128 75454
rect 507808 75134 508128 75218
rect 507808 74898 507850 75134
rect 508086 74898 508128 75134
rect 507808 74866 508128 74898
rect 538528 75454 538848 75486
rect 538528 75218 538570 75454
rect 538806 75218 538848 75454
rect 538528 75134 538848 75218
rect 538528 74898 538570 75134
rect 538806 74898 538848 75134
rect 538528 74866 538848 74898
rect 62368 57454 62688 57486
rect 62368 57218 62410 57454
rect 62646 57218 62688 57454
rect 62368 57134 62688 57218
rect 62368 56898 62410 57134
rect 62646 56898 62688 57134
rect 62368 56866 62688 56898
rect 93088 57454 93408 57486
rect 93088 57218 93130 57454
rect 93366 57218 93408 57454
rect 93088 57134 93408 57218
rect 93088 56898 93130 57134
rect 93366 56898 93408 57134
rect 93088 56866 93408 56898
rect 123808 57454 124128 57486
rect 123808 57218 123850 57454
rect 124086 57218 124128 57454
rect 123808 57134 124128 57218
rect 123808 56898 123850 57134
rect 124086 56898 124128 57134
rect 123808 56866 124128 56898
rect 154528 57454 154848 57486
rect 154528 57218 154570 57454
rect 154806 57218 154848 57454
rect 154528 57134 154848 57218
rect 154528 56898 154570 57134
rect 154806 56898 154848 57134
rect 154528 56866 154848 56898
rect 185248 57454 185568 57486
rect 185248 57218 185290 57454
rect 185526 57218 185568 57454
rect 185248 57134 185568 57218
rect 185248 56898 185290 57134
rect 185526 56898 185568 57134
rect 185248 56866 185568 56898
rect 215968 57454 216288 57486
rect 215968 57218 216010 57454
rect 216246 57218 216288 57454
rect 215968 57134 216288 57218
rect 215968 56898 216010 57134
rect 216246 56898 216288 57134
rect 215968 56866 216288 56898
rect 246688 57454 247008 57486
rect 246688 57218 246730 57454
rect 246966 57218 247008 57454
rect 246688 57134 247008 57218
rect 246688 56898 246730 57134
rect 246966 56898 247008 57134
rect 246688 56866 247008 56898
rect 277408 57454 277728 57486
rect 277408 57218 277450 57454
rect 277686 57218 277728 57454
rect 277408 57134 277728 57218
rect 277408 56898 277450 57134
rect 277686 56898 277728 57134
rect 277408 56866 277728 56898
rect 308128 57454 308448 57486
rect 308128 57218 308170 57454
rect 308406 57218 308448 57454
rect 308128 57134 308448 57218
rect 308128 56898 308170 57134
rect 308406 56898 308448 57134
rect 308128 56866 308448 56898
rect 338848 57454 339168 57486
rect 338848 57218 338890 57454
rect 339126 57218 339168 57454
rect 338848 57134 339168 57218
rect 338848 56898 338890 57134
rect 339126 56898 339168 57134
rect 338848 56866 339168 56898
rect 369568 57454 369888 57486
rect 369568 57218 369610 57454
rect 369846 57218 369888 57454
rect 369568 57134 369888 57218
rect 369568 56898 369610 57134
rect 369846 56898 369888 57134
rect 369568 56866 369888 56898
rect 400288 57454 400608 57486
rect 400288 57218 400330 57454
rect 400566 57218 400608 57454
rect 400288 57134 400608 57218
rect 400288 56898 400330 57134
rect 400566 56898 400608 57134
rect 400288 56866 400608 56898
rect 431008 57454 431328 57486
rect 431008 57218 431050 57454
rect 431286 57218 431328 57454
rect 431008 57134 431328 57218
rect 431008 56898 431050 57134
rect 431286 56898 431328 57134
rect 431008 56866 431328 56898
rect 461728 57454 462048 57486
rect 461728 57218 461770 57454
rect 462006 57218 462048 57454
rect 461728 57134 462048 57218
rect 461728 56898 461770 57134
rect 462006 56898 462048 57134
rect 461728 56866 462048 56898
rect 492448 57454 492768 57486
rect 492448 57218 492490 57454
rect 492726 57218 492768 57454
rect 492448 57134 492768 57218
rect 492448 56898 492490 57134
rect 492726 56898 492768 57134
rect 492448 56866 492768 56898
rect 523168 57454 523488 57486
rect 523168 57218 523210 57454
rect 523446 57218 523488 57454
rect 523168 57134 523488 57218
rect 523168 56898 523210 57134
rect 523446 56898 523488 57134
rect 523168 56866 523488 56898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 43174 42134 51000
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 46894 45854 51000
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 50614 49574 51000
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 51000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 51000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 51000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 51000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 51000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 51000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 51000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 51000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 51000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 51000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 51000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 51000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 51000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 51000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 51000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 51000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 51000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 51000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 51000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 51000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 51000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 51000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 51000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 51000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 51000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 51000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 51000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 51000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 51000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 51000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 51000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 51000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 51000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 51000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 51000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 51000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 51000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 51000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 51000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 51000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 51000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 51000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 51000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 51000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 51000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 51000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 51000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 51000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 51000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 51000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 51000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 51000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 51000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 51000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 51000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 51000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 51000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 51000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 51000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 51000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 51000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 51000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 51000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 51000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 51000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 51000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 51000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 51000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 51000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 51000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 51000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 51000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 51000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 51000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 51000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 51000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 51000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 51000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 51000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 51000
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 51000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 51000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 51000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 51000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 51000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 51000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 51000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 51000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 51000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 51000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 51000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 51000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 51000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 51000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 51000
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 51000
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 51000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 51000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 51000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 51000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 51000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 51000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 51000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 51000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 51000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 51000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 28894 531854 51000
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 32614 535574 51000
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 39454 542414 51000
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 43174 546134 51000
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 47050 651218 47286 651454
rect 47050 650898 47286 651134
rect 77770 651218 78006 651454
rect 77770 650898 78006 651134
rect 108490 651218 108726 651454
rect 108490 650898 108726 651134
rect 139210 651218 139446 651454
rect 139210 650898 139446 651134
rect 169930 651218 170166 651454
rect 169930 650898 170166 651134
rect 200650 651218 200886 651454
rect 200650 650898 200886 651134
rect 231370 651218 231606 651454
rect 231370 650898 231606 651134
rect 262090 651218 262326 651454
rect 262090 650898 262326 651134
rect 292810 651218 293046 651454
rect 292810 650898 293046 651134
rect 323530 651218 323766 651454
rect 323530 650898 323766 651134
rect 354250 651218 354486 651454
rect 354250 650898 354486 651134
rect 384970 651218 385206 651454
rect 384970 650898 385206 651134
rect 415690 651218 415926 651454
rect 415690 650898 415926 651134
rect 446410 651218 446646 651454
rect 446410 650898 446646 651134
rect 477130 651218 477366 651454
rect 477130 650898 477366 651134
rect 507850 651218 508086 651454
rect 507850 650898 508086 651134
rect 538570 651218 538806 651454
rect 538570 650898 538806 651134
rect 62410 633218 62646 633454
rect 62410 632898 62646 633134
rect 93130 633218 93366 633454
rect 93130 632898 93366 633134
rect 123850 633218 124086 633454
rect 123850 632898 124086 633134
rect 154570 633218 154806 633454
rect 154570 632898 154806 633134
rect 185290 633218 185526 633454
rect 185290 632898 185526 633134
rect 216010 633218 216246 633454
rect 216010 632898 216246 633134
rect 246730 633218 246966 633454
rect 246730 632898 246966 633134
rect 277450 633218 277686 633454
rect 277450 632898 277686 633134
rect 308170 633218 308406 633454
rect 308170 632898 308406 633134
rect 338890 633218 339126 633454
rect 338890 632898 339126 633134
rect 369610 633218 369846 633454
rect 369610 632898 369846 633134
rect 400330 633218 400566 633454
rect 400330 632898 400566 633134
rect 431050 633218 431286 633454
rect 431050 632898 431286 633134
rect 461770 633218 462006 633454
rect 461770 632898 462006 633134
rect 492490 633218 492726 633454
rect 492490 632898 492726 633134
rect 523210 633218 523446 633454
rect 523210 632898 523446 633134
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 47050 615218 47286 615454
rect 47050 614898 47286 615134
rect 77770 615218 78006 615454
rect 77770 614898 78006 615134
rect 108490 615218 108726 615454
rect 108490 614898 108726 615134
rect 139210 615218 139446 615454
rect 139210 614898 139446 615134
rect 169930 615218 170166 615454
rect 169930 614898 170166 615134
rect 200650 615218 200886 615454
rect 200650 614898 200886 615134
rect 231370 615218 231606 615454
rect 231370 614898 231606 615134
rect 262090 615218 262326 615454
rect 262090 614898 262326 615134
rect 292810 615218 293046 615454
rect 292810 614898 293046 615134
rect 323530 615218 323766 615454
rect 323530 614898 323766 615134
rect 354250 615218 354486 615454
rect 354250 614898 354486 615134
rect 384970 615218 385206 615454
rect 384970 614898 385206 615134
rect 415690 615218 415926 615454
rect 415690 614898 415926 615134
rect 446410 615218 446646 615454
rect 446410 614898 446646 615134
rect 477130 615218 477366 615454
rect 477130 614898 477366 615134
rect 507850 615218 508086 615454
rect 507850 614898 508086 615134
rect 538570 615218 538806 615454
rect 538570 614898 538806 615134
rect 62410 597218 62646 597454
rect 62410 596898 62646 597134
rect 93130 597218 93366 597454
rect 93130 596898 93366 597134
rect 123850 597218 124086 597454
rect 123850 596898 124086 597134
rect 154570 597218 154806 597454
rect 154570 596898 154806 597134
rect 185290 597218 185526 597454
rect 185290 596898 185526 597134
rect 216010 597218 216246 597454
rect 216010 596898 216246 597134
rect 246730 597218 246966 597454
rect 246730 596898 246966 597134
rect 277450 597218 277686 597454
rect 277450 596898 277686 597134
rect 308170 597218 308406 597454
rect 308170 596898 308406 597134
rect 338890 597218 339126 597454
rect 338890 596898 339126 597134
rect 369610 597218 369846 597454
rect 369610 596898 369846 597134
rect 400330 597218 400566 597454
rect 400330 596898 400566 597134
rect 431050 597218 431286 597454
rect 431050 596898 431286 597134
rect 461770 597218 462006 597454
rect 461770 596898 462006 597134
rect 492490 597218 492726 597454
rect 492490 596898 492726 597134
rect 523210 597218 523446 597454
rect 523210 596898 523446 597134
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 47050 579218 47286 579454
rect 47050 578898 47286 579134
rect 77770 579218 78006 579454
rect 77770 578898 78006 579134
rect 108490 579218 108726 579454
rect 108490 578898 108726 579134
rect 139210 579218 139446 579454
rect 139210 578898 139446 579134
rect 169930 579218 170166 579454
rect 169930 578898 170166 579134
rect 200650 579218 200886 579454
rect 200650 578898 200886 579134
rect 231370 579218 231606 579454
rect 231370 578898 231606 579134
rect 262090 579218 262326 579454
rect 262090 578898 262326 579134
rect 292810 579218 293046 579454
rect 292810 578898 293046 579134
rect 323530 579218 323766 579454
rect 323530 578898 323766 579134
rect 354250 579218 354486 579454
rect 354250 578898 354486 579134
rect 384970 579218 385206 579454
rect 384970 578898 385206 579134
rect 415690 579218 415926 579454
rect 415690 578898 415926 579134
rect 446410 579218 446646 579454
rect 446410 578898 446646 579134
rect 477130 579218 477366 579454
rect 477130 578898 477366 579134
rect 507850 579218 508086 579454
rect 507850 578898 508086 579134
rect 538570 579218 538806 579454
rect 538570 578898 538806 579134
rect 62410 561218 62646 561454
rect 62410 560898 62646 561134
rect 93130 561218 93366 561454
rect 93130 560898 93366 561134
rect 123850 561218 124086 561454
rect 123850 560898 124086 561134
rect 154570 561218 154806 561454
rect 154570 560898 154806 561134
rect 185290 561218 185526 561454
rect 185290 560898 185526 561134
rect 216010 561218 216246 561454
rect 216010 560898 216246 561134
rect 246730 561218 246966 561454
rect 246730 560898 246966 561134
rect 277450 561218 277686 561454
rect 277450 560898 277686 561134
rect 308170 561218 308406 561454
rect 308170 560898 308406 561134
rect 338890 561218 339126 561454
rect 338890 560898 339126 561134
rect 369610 561218 369846 561454
rect 369610 560898 369846 561134
rect 400330 561218 400566 561454
rect 400330 560898 400566 561134
rect 431050 561218 431286 561454
rect 431050 560898 431286 561134
rect 461770 561218 462006 561454
rect 461770 560898 462006 561134
rect 492490 561218 492726 561454
rect 492490 560898 492726 561134
rect 523210 561218 523446 561454
rect 523210 560898 523446 561134
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 47050 543218 47286 543454
rect 47050 542898 47286 543134
rect 77770 543218 78006 543454
rect 77770 542898 78006 543134
rect 108490 543218 108726 543454
rect 108490 542898 108726 543134
rect 139210 543218 139446 543454
rect 139210 542898 139446 543134
rect 169930 543218 170166 543454
rect 169930 542898 170166 543134
rect 200650 543218 200886 543454
rect 200650 542898 200886 543134
rect 231370 543218 231606 543454
rect 231370 542898 231606 543134
rect 262090 543218 262326 543454
rect 262090 542898 262326 543134
rect 292810 543218 293046 543454
rect 292810 542898 293046 543134
rect 323530 543218 323766 543454
rect 323530 542898 323766 543134
rect 354250 543218 354486 543454
rect 354250 542898 354486 543134
rect 384970 543218 385206 543454
rect 384970 542898 385206 543134
rect 415690 543218 415926 543454
rect 415690 542898 415926 543134
rect 446410 543218 446646 543454
rect 446410 542898 446646 543134
rect 477130 543218 477366 543454
rect 477130 542898 477366 543134
rect 507850 543218 508086 543454
rect 507850 542898 508086 543134
rect 538570 543218 538806 543454
rect 538570 542898 538806 543134
rect 62410 525218 62646 525454
rect 62410 524898 62646 525134
rect 93130 525218 93366 525454
rect 93130 524898 93366 525134
rect 123850 525218 124086 525454
rect 123850 524898 124086 525134
rect 154570 525218 154806 525454
rect 154570 524898 154806 525134
rect 185290 525218 185526 525454
rect 185290 524898 185526 525134
rect 216010 525218 216246 525454
rect 216010 524898 216246 525134
rect 246730 525218 246966 525454
rect 246730 524898 246966 525134
rect 277450 525218 277686 525454
rect 277450 524898 277686 525134
rect 308170 525218 308406 525454
rect 308170 524898 308406 525134
rect 338890 525218 339126 525454
rect 338890 524898 339126 525134
rect 369610 525218 369846 525454
rect 369610 524898 369846 525134
rect 400330 525218 400566 525454
rect 400330 524898 400566 525134
rect 431050 525218 431286 525454
rect 431050 524898 431286 525134
rect 461770 525218 462006 525454
rect 461770 524898 462006 525134
rect 492490 525218 492726 525454
rect 492490 524898 492726 525134
rect 523210 525218 523446 525454
rect 523210 524898 523446 525134
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 47050 507218 47286 507454
rect 47050 506898 47286 507134
rect 77770 507218 78006 507454
rect 77770 506898 78006 507134
rect 108490 507218 108726 507454
rect 108490 506898 108726 507134
rect 139210 507218 139446 507454
rect 139210 506898 139446 507134
rect 169930 507218 170166 507454
rect 169930 506898 170166 507134
rect 200650 507218 200886 507454
rect 200650 506898 200886 507134
rect 231370 507218 231606 507454
rect 231370 506898 231606 507134
rect 262090 507218 262326 507454
rect 262090 506898 262326 507134
rect 292810 507218 293046 507454
rect 292810 506898 293046 507134
rect 323530 507218 323766 507454
rect 323530 506898 323766 507134
rect 354250 507218 354486 507454
rect 354250 506898 354486 507134
rect 384970 507218 385206 507454
rect 384970 506898 385206 507134
rect 415690 507218 415926 507454
rect 415690 506898 415926 507134
rect 446410 507218 446646 507454
rect 446410 506898 446646 507134
rect 477130 507218 477366 507454
rect 477130 506898 477366 507134
rect 507850 507218 508086 507454
rect 507850 506898 508086 507134
rect 538570 507218 538806 507454
rect 538570 506898 538806 507134
rect 62410 489218 62646 489454
rect 62410 488898 62646 489134
rect 93130 489218 93366 489454
rect 93130 488898 93366 489134
rect 123850 489218 124086 489454
rect 123850 488898 124086 489134
rect 154570 489218 154806 489454
rect 154570 488898 154806 489134
rect 185290 489218 185526 489454
rect 185290 488898 185526 489134
rect 216010 489218 216246 489454
rect 216010 488898 216246 489134
rect 246730 489218 246966 489454
rect 246730 488898 246966 489134
rect 277450 489218 277686 489454
rect 277450 488898 277686 489134
rect 308170 489218 308406 489454
rect 308170 488898 308406 489134
rect 338890 489218 339126 489454
rect 338890 488898 339126 489134
rect 369610 489218 369846 489454
rect 369610 488898 369846 489134
rect 400330 489218 400566 489454
rect 400330 488898 400566 489134
rect 431050 489218 431286 489454
rect 431050 488898 431286 489134
rect 461770 489218 462006 489454
rect 461770 488898 462006 489134
rect 492490 489218 492726 489454
rect 492490 488898 492726 489134
rect 523210 489218 523446 489454
rect 523210 488898 523446 489134
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 47050 471218 47286 471454
rect 47050 470898 47286 471134
rect 77770 471218 78006 471454
rect 77770 470898 78006 471134
rect 108490 471218 108726 471454
rect 108490 470898 108726 471134
rect 139210 471218 139446 471454
rect 139210 470898 139446 471134
rect 169930 471218 170166 471454
rect 169930 470898 170166 471134
rect 200650 471218 200886 471454
rect 200650 470898 200886 471134
rect 231370 471218 231606 471454
rect 231370 470898 231606 471134
rect 262090 471218 262326 471454
rect 262090 470898 262326 471134
rect 292810 471218 293046 471454
rect 292810 470898 293046 471134
rect 323530 471218 323766 471454
rect 323530 470898 323766 471134
rect 354250 471218 354486 471454
rect 354250 470898 354486 471134
rect 384970 471218 385206 471454
rect 384970 470898 385206 471134
rect 415690 471218 415926 471454
rect 415690 470898 415926 471134
rect 446410 471218 446646 471454
rect 446410 470898 446646 471134
rect 477130 471218 477366 471454
rect 477130 470898 477366 471134
rect 507850 471218 508086 471454
rect 507850 470898 508086 471134
rect 538570 471218 538806 471454
rect 538570 470898 538806 471134
rect 62410 453218 62646 453454
rect 62410 452898 62646 453134
rect 93130 453218 93366 453454
rect 93130 452898 93366 453134
rect 123850 453218 124086 453454
rect 123850 452898 124086 453134
rect 154570 453218 154806 453454
rect 154570 452898 154806 453134
rect 185290 453218 185526 453454
rect 185290 452898 185526 453134
rect 216010 453218 216246 453454
rect 216010 452898 216246 453134
rect 246730 453218 246966 453454
rect 246730 452898 246966 453134
rect 277450 453218 277686 453454
rect 277450 452898 277686 453134
rect 308170 453218 308406 453454
rect 308170 452898 308406 453134
rect 338890 453218 339126 453454
rect 338890 452898 339126 453134
rect 369610 453218 369846 453454
rect 369610 452898 369846 453134
rect 400330 453218 400566 453454
rect 400330 452898 400566 453134
rect 431050 453218 431286 453454
rect 431050 452898 431286 453134
rect 461770 453218 462006 453454
rect 461770 452898 462006 453134
rect 492490 453218 492726 453454
rect 492490 452898 492726 453134
rect 523210 453218 523446 453454
rect 523210 452898 523446 453134
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 47050 435218 47286 435454
rect 47050 434898 47286 435134
rect 77770 435218 78006 435454
rect 77770 434898 78006 435134
rect 108490 435218 108726 435454
rect 108490 434898 108726 435134
rect 139210 435218 139446 435454
rect 139210 434898 139446 435134
rect 169930 435218 170166 435454
rect 169930 434898 170166 435134
rect 200650 435218 200886 435454
rect 200650 434898 200886 435134
rect 231370 435218 231606 435454
rect 231370 434898 231606 435134
rect 262090 435218 262326 435454
rect 262090 434898 262326 435134
rect 292810 435218 293046 435454
rect 292810 434898 293046 435134
rect 323530 435218 323766 435454
rect 323530 434898 323766 435134
rect 354250 435218 354486 435454
rect 354250 434898 354486 435134
rect 384970 435218 385206 435454
rect 384970 434898 385206 435134
rect 415690 435218 415926 435454
rect 415690 434898 415926 435134
rect 446410 435218 446646 435454
rect 446410 434898 446646 435134
rect 477130 435218 477366 435454
rect 477130 434898 477366 435134
rect 507850 435218 508086 435454
rect 507850 434898 508086 435134
rect 538570 435218 538806 435454
rect 538570 434898 538806 435134
rect 62410 417218 62646 417454
rect 62410 416898 62646 417134
rect 93130 417218 93366 417454
rect 93130 416898 93366 417134
rect 123850 417218 124086 417454
rect 123850 416898 124086 417134
rect 154570 417218 154806 417454
rect 154570 416898 154806 417134
rect 185290 417218 185526 417454
rect 185290 416898 185526 417134
rect 216010 417218 216246 417454
rect 216010 416898 216246 417134
rect 246730 417218 246966 417454
rect 246730 416898 246966 417134
rect 277450 417218 277686 417454
rect 277450 416898 277686 417134
rect 308170 417218 308406 417454
rect 308170 416898 308406 417134
rect 338890 417218 339126 417454
rect 338890 416898 339126 417134
rect 369610 417218 369846 417454
rect 369610 416898 369846 417134
rect 400330 417218 400566 417454
rect 400330 416898 400566 417134
rect 431050 417218 431286 417454
rect 431050 416898 431286 417134
rect 461770 417218 462006 417454
rect 461770 416898 462006 417134
rect 492490 417218 492726 417454
rect 492490 416898 492726 417134
rect 523210 417218 523446 417454
rect 523210 416898 523446 417134
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 47050 399218 47286 399454
rect 47050 398898 47286 399134
rect 77770 399218 78006 399454
rect 77770 398898 78006 399134
rect 108490 399218 108726 399454
rect 108490 398898 108726 399134
rect 139210 399218 139446 399454
rect 139210 398898 139446 399134
rect 169930 399218 170166 399454
rect 169930 398898 170166 399134
rect 200650 399218 200886 399454
rect 200650 398898 200886 399134
rect 231370 399218 231606 399454
rect 231370 398898 231606 399134
rect 262090 399218 262326 399454
rect 262090 398898 262326 399134
rect 292810 399218 293046 399454
rect 292810 398898 293046 399134
rect 323530 399218 323766 399454
rect 323530 398898 323766 399134
rect 354250 399218 354486 399454
rect 354250 398898 354486 399134
rect 384970 399218 385206 399454
rect 384970 398898 385206 399134
rect 415690 399218 415926 399454
rect 415690 398898 415926 399134
rect 446410 399218 446646 399454
rect 446410 398898 446646 399134
rect 477130 399218 477366 399454
rect 477130 398898 477366 399134
rect 507850 399218 508086 399454
rect 507850 398898 508086 399134
rect 538570 399218 538806 399454
rect 538570 398898 538806 399134
rect 62410 381218 62646 381454
rect 62410 380898 62646 381134
rect 93130 381218 93366 381454
rect 93130 380898 93366 381134
rect 123850 381218 124086 381454
rect 123850 380898 124086 381134
rect 154570 381218 154806 381454
rect 154570 380898 154806 381134
rect 185290 381218 185526 381454
rect 185290 380898 185526 381134
rect 216010 381218 216246 381454
rect 216010 380898 216246 381134
rect 246730 381218 246966 381454
rect 246730 380898 246966 381134
rect 277450 381218 277686 381454
rect 277450 380898 277686 381134
rect 308170 381218 308406 381454
rect 308170 380898 308406 381134
rect 338890 381218 339126 381454
rect 338890 380898 339126 381134
rect 369610 381218 369846 381454
rect 369610 380898 369846 381134
rect 400330 381218 400566 381454
rect 400330 380898 400566 381134
rect 431050 381218 431286 381454
rect 431050 380898 431286 381134
rect 461770 381218 462006 381454
rect 461770 380898 462006 381134
rect 492490 381218 492726 381454
rect 492490 380898 492726 381134
rect 523210 381218 523446 381454
rect 523210 380898 523446 381134
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 47050 363218 47286 363454
rect 47050 362898 47286 363134
rect 77770 363218 78006 363454
rect 77770 362898 78006 363134
rect 108490 363218 108726 363454
rect 108490 362898 108726 363134
rect 139210 363218 139446 363454
rect 139210 362898 139446 363134
rect 169930 363218 170166 363454
rect 169930 362898 170166 363134
rect 200650 363218 200886 363454
rect 200650 362898 200886 363134
rect 231370 363218 231606 363454
rect 231370 362898 231606 363134
rect 262090 363218 262326 363454
rect 262090 362898 262326 363134
rect 292810 363218 293046 363454
rect 292810 362898 293046 363134
rect 323530 363218 323766 363454
rect 323530 362898 323766 363134
rect 354250 363218 354486 363454
rect 354250 362898 354486 363134
rect 384970 363218 385206 363454
rect 384970 362898 385206 363134
rect 415690 363218 415926 363454
rect 415690 362898 415926 363134
rect 446410 363218 446646 363454
rect 446410 362898 446646 363134
rect 477130 363218 477366 363454
rect 477130 362898 477366 363134
rect 507850 363218 508086 363454
rect 507850 362898 508086 363134
rect 538570 363218 538806 363454
rect 538570 362898 538806 363134
rect 62410 345218 62646 345454
rect 62410 344898 62646 345134
rect 93130 345218 93366 345454
rect 93130 344898 93366 345134
rect 123850 345218 124086 345454
rect 123850 344898 124086 345134
rect 154570 345218 154806 345454
rect 154570 344898 154806 345134
rect 185290 345218 185526 345454
rect 185290 344898 185526 345134
rect 216010 345218 216246 345454
rect 216010 344898 216246 345134
rect 246730 345218 246966 345454
rect 246730 344898 246966 345134
rect 277450 345218 277686 345454
rect 277450 344898 277686 345134
rect 308170 345218 308406 345454
rect 308170 344898 308406 345134
rect 338890 345218 339126 345454
rect 338890 344898 339126 345134
rect 369610 345218 369846 345454
rect 369610 344898 369846 345134
rect 400330 345218 400566 345454
rect 400330 344898 400566 345134
rect 431050 345218 431286 345454
rect 431050 344898 431286 345134
rect 461770 345218 462006 345454
rect 461770 344898 462006 345134
rect 492490 345218 492726 345454
rect 492490 344898 492726 345134
rect 523210 345218 523446 345454
rect 523210 344898 523446 345134
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 47050 327218 47286 327454
rect 47050 326898 47286 327134
rect 77770 327218 78006 327454
rect 77770 326898 78006 327134
rect 108490 327218 108726 327454
rect 108490 326898 108726 327134
rect 139210 327218 139446 327454
rect 139210 326898 139446 327134
rect 169930 327218 170166 327454
rect 169930 326898 170166 327134
rect 200650 327218 200886 327454
rect 200650 326898 200886 327134
rect 231370 327218 231606 327454
rect 231370 326898 231606 327134
rect 262090 327218 262326 327454
rect 262090 326898 262326 327134
rect 292810 327218 293046 327454
rect 292810 326898 293046 327134
rect 323530 327218 323766 327454
rect 323530 326898 323766 327134
rect 354250 327218 354486 327454
rect 354250 326898 354486 327134
rect 384970 327218 385206 327454
rect 384970 326898 385206 327134
rect 415690 327218 415926 327454
rect 415690 326898 415926 327134
rect 446410 327218 446646 327454
rect 446410 326898 446646 327134
rect 477130 327218 477366 327454
rect 477130 326898 477366 327134
rect 507850 327218 508086 327454
rect 507850 326898 508086 327134
rect 538570 327218 538806 327454
rect 538570 326898 538806 327134
rect 62410 309218 62646 309454
rect 62410 308898 62646 309134
rect 93130 309218 93366 309454
rect 93130 308898 93366 309134
rect 123850 309218 124086 309454
rect 123850 308898 124086 309134
rect 154570 309218 154806 309454
rect 154570 308898 154806 309134
rect 185290 309218 185526 309454
rect 185290 308898 185526 309134
rect 216010 309218 216246 309454
rect 216010 308898 216246 309134
rect 246730 309218 246966 309454
rect 246730 308898 246966 309134
rect 277450 309218 277686 309454
rect 277450 308898 277686 309134
rect 308170 309218 308406 309454
rect 308170 308898 308406 309134
rect 338890 309218 339126 309454
rect 338890 308898 339126 309134
rect 369610 309218 369846 309454
rect 369610 308898 369846 309134
rect 400330 309218 400566 309454
rect 400330 308898 400566 309134
rect 431050 309218 431286 309454
rect 431050 308898 431286 309134
rect 461770 309218 462006 309454
rect 461770 308898 462006 309134
rect 492490 309218 492726 309454
rect 492490 308898 492726 309134
rect 523210 309218 523446 309454
rect 523210 308898 523446 309134
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 47050 291218 47286 291454
rect 47050 290898 47286 291134
rect 77770 291218 78006 291454
rect 77770 290898 78006 291134
rect 108490 291218 108726 291454
rect 108490 290898 108726 291134
rect 139210 291218 139446 291454
rect 139210 290898 139446 291134
rect 169930 291218 170166 291454
rect 169930 290898 170166 291134
rect 200650 291218 200886 291454
rect 200650 290898 200886 291134
rect 231370 291218 231606 291454
rect 231370 290898 231606 291134
rect 262090 291218 262326 291454
rect 262090 290898 262326 291134
rect 292810 291218 293046 291454
rect 292810 290898 293046 291134
rect 323530 291218 323766 291454
rect 323530 290898 323766 291134
rect 354250 291218 354486 291454
rect 354250 290898 354486 291134
rect 384970 291218 385206 291454
rect 384970 290898 385206 291134
rect 415690 291218 415926 291454
rect 415690 290898 415926 291134
rect 446410 291218 446646 291454
rect 446410 290898 446646 291134
rect 477130 291218 477366 291454
rect 477130 290898 477366 291134
rect 507850 291218 508086 291454
rect 507850 290898 508086 291134
rect 538570 291218 538806 291454
rect 538570 290898 538806 291134
rect 62410 273218 62646 273454
rect 62410 272898 62646 273134
rect 93130 273218 93366 273454
rect 93130 272898 93366 273134
rect 123850 273218 124086 273454
rect 123850 272898 124086 273134
rect 154570 273218 154806 273454
rect 154570 272898 154806 273134
rect 185290 273218 185526 273454
rect 185290 272898 185526 273134
rect 216010 273218 216246 273454
rect 216010 272898 216246 273134
rect 246730 273218 246966 273454
rect 246730 272898 246966 273134
rect 277450 273218 277686 273454
rect 277450 272898 277686 273134
rect 308170 273218 308406 273454
rect 308170 272898 308406 273134
rect 338890 273218 339126 273454
rect 338890 272898 339126 273134
rect 369610 273218 369846 273454
rect 369610 272898 369846 273134
rect 400330 273218 400566 273454
rect 400330 272898 400566 273134
rect 431050 273218 431286 273454
rect 431050 272898 431286 273134
rect 461770 273218 462006 273454
rect 461770 272898 462006 273134
rect 492490 273218 492726 273454
rect 492490 272898 492726 273134
rect 523210 273218 523446 273454
rect 523210 272898 523446 273134
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 47050 255218 47286 255454
rect 47050 254898 47286 255134
rect 77770 255218 78006 255454
rect 77770 254898 78006 255134
rect 108490 255218 108726 255454
rect 108490 254898 108726 255134
rect 139210 255218 139446 255454
rect 139210 254898 139446 255134
rect 169930 255218 170166 255454
rect 169930 254898 170166 255134
rect 200650 255218 200886 255454
rect 200650 254898 200886 255134
rect 231370 255218 231606 255454
rect 231370 254898 231606 255134
rect 262090 255218 262326 255454
rect 262090 254898 262326 255134
rect 292810 255218 293046 255454
rect 292810 254898 293046 255134
rect 323530 255218 323766 255454
rect 323530 254898 323766 255134
rect 354250 255218 354486 255454
rect 354250 254898 354486 255134
rect 384970 255218 385206 255454
rect 384970 254898 385206 255134
rect 415690 255218 415926 255454
rect 415690 254898 415926 255134
rect 446410 255218 446646 255454
rect 446410 254898 446646 255134
rect 477130 255218 477366 255454
rect 477130 254898 477366 255134
rect 507850 255218 508086 255454
rect 507850 254898 508086 255134
rect 538570 255218 538806 255454
rect 538570 254898 538806 255134
rect 62410 237218 62646 237454
rect 62410 236898 62646 237134
rect 93130 237218 93366 237454
rect 93130 236898 93366 237134
rect 123850 237218 124086 237454
rect 123850 236898 124086 237134
rect 154570 237218 154806 237454
rect 154570 236898 154806 237134
rect 185290 237218 185526 237454
rect 185290 236898 185526 237134
rect 216010 237218 216246 237454
rect 216010 236898 216246 237134
rect 246730 237218 246966 237454
rect 246730 236898 246966 237134
rect 277450 237218 277686 237454
rect 277450 236898 277686 237134
rect 308170 237218 308406 237454
rect 308170 236898 308406 237134
rect 338890 237218 339126 237454
rect 338890 236898 339126 237134
rect 369610 237218 369846 237454
rect 369610 236898 369846 237134
rect 400330 237218 400566 237454
rect 400330 236898 400566 237134
rect 431050 237218 431286 237454
rect 431050 236898 431286 237134
rect 461770 237218 462006 237454
rect 461770 236898 462006 237134
rect 492490 237218 492726 237454
rect 492490 236898 492726 237134
rect 523210 237218 523446 237454
rect 523210 236898 523446 237134
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 47050 219218 47286 219454
rect 47050 218898 47286 219134
rect 77770 219218 78006 219454
rect 77770 218898 78006 219134
rect 108490 219218 108726 219454
rect 108490 218898 108726 219134
rect 139210 219218 139446 219454
rect 139210 218898 139446 219134
rect 169930 219218 170166 219454
rect 169930 218898 170166 219134
rect 200650 219218 200886 219454
rect 200650 218898 200886 219134
rect 231370 219218 231606 219454
rect 231370 218898 231606 219134
rect 262090 219218 262326 219454
rect 262090 218898 262326 219134
rect 292810 219218 293046 219454
rect 292810 218898 293046 219134
rect 323530 219218 323766 219454
rect 323530 218898 323766 219134
rect 354250 219218 354486 219454
rect 354250 218898 354486 219134
rect 384970 219218 385206 219454
rect 384970 218898 385206 219134
rect 415690 219218 415926 219454
rect 415690 218898 415926 219134
rect 446410 219218 446646 219454
rect 446410 218898 446646 219134
rect 477130 219218 477366 219454
rect 477130 218898 477366 219134
rect 507850 219218 508086 219454
rect 507850 218898 508086 219134
rect 538570 219218 538806 219454
rect 538570 218898 538806 219134
rect 62410 201218 62646 201454
rect 62410 200898 62646 201134
rect 93130 201218 93366 201454
rect 93130 200898 93366 201134
rect 123850 201218 124086 201454
rect 123850 200898 124086 201134
rect 154570 201218 154806 201454
rect 154570 200898 154806 201134
rect 185290 201218 185526 201454
rect 185290 200898 185526 201134
rect 216010 201218 216246 201454
rect 216010 200898 216246 201134
rect 246730 201218 246966 201454
rect 246730 200898 246966 201134
rect 277450 201218 277686 201454
rect 277450 200898 277686 201134
rect 308170 201218 308406 201454
rect 308170 200898 308406 201134
rect 338890 201218 339126 201454
rect 338890 200898 339126 201134
rect 369610 201218 369846 201454
rect 369610 200898 369846 201134
rect 400330 201218 400566 201454
rect 400330 200898 400566 201134
rect 431050 201218 431286 201454
rect 431050 200898 431286 201134
rect 461770 201218 462006 201454
rect 461770 200898 462006 201134
rect 492490 201218 492726 201454
rect 492490 200898 492726 201134
rect 523210 201218 523446 201454
rect 523210 200898 523446 201134
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 47050 183218 47286 183454
rect 47050 182898 47286 183134
rect 77770 183218 78006 183454
rect 77770 182898 78006 183134
rect 108490 183218 108726 183454
rect 108490 182898 108726 183134
rect 139210 183218 139446 183454
rect 139210 182898 139446 183134
rect 169930 183218 170166 183454
rect 169930 182898 170166 183134
rect 200650 183218 200886 183454
rect 200650 182898 200886 183134
rect 231370 183218 231606 183454
rect 231370 182898 231606 183134
rect 262090 183218 262326 183454
rect 262090 182898 262326 183134
rect 292810 183218 293046 183454
rect 292810 182898 293046 183134
rect 323530 183218 323766 183454
rect 323530 182898 323766 183134
rect 354250 183218 354486 183454
rect 354250 182898 354486 183134
rect 384970 183218 385206 183454
rect 384970 182898 385206 183134
rect 415690 183218 415926 183454
rect 415690 182898 415926 183134
rect 446410 183218 446646 183454
rect 446410 182898 446646 183134
rect 477130 183218 477366 183454
rect 477130 182898 477366 183134
rect 507850 183218 508086 183454
rect 507850 182898 508086 183134
rect 538570 183218 538806 183454
rect 538570 182898 538806 183134
rect 62410 165218 62646 165454
rect 62410 164898 62646 165134
rect 93130 165218 93366 165454
rect 93130 164898 93366 165134
rect 123850 165218 124086 165454
rect 123850 164898 124086 165134
rect 154570 165218 154806 165454
rect 154570 164898 154806 165134
rect 185290 165218 185526 165454
rect 185290 164898 185526 165134
rect 216010 165218 216246 165454
rect 216010 164898 216246 165134
rect 246730 165218 246966 165454
rect 246730 164898 246966 165134
rect 277450 165218 277686 165454
rect 277450 164898 277686 165134
rect 308170 165218 308406 165454
rect 308170 164898 308406 165134
rect 338890 165218 339126 165454
rect 338890 164898 339126 165134
rect 369610 165218 369846 165454
rect 369610 164898 369846 165134
rect 400330 165218 400566 165454
rect 400330 164898 400566 165134
rect 431050 165218 431286 165454
rect 431050 164898 431286 165134
rect 461770 165218 462006 165454
rect 461770 164898 462006 165134
rect 492490 165218 492726 165454
rect 492490 164898 492726 165134
rect 523210 165218 523446 165454
rect 523210 164898 523446 165134
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 47050 147218 47286 147454
rect 47050 146898 47286 147134
rect 77770 147218 78006 147454
rect 77770 146898 78006 147134
rect 108490 147218 108726 147454
rect 108490 146898 108726 147134
rect 139210 147218 139446 147454
rect 139210 146898 139446 147134
rect 169930 147218 170166 147454
rect 169930 146898 170166 147134
rect 200650 147218 200886 147454
rect 200650 146898 200886 147134
rect 231370 147218 231606 147454
rect 231370 146898 231606 147134
rect 262090 147218 262326 147454
rect 262090 146898 262326 147134
rect 292810 147218 293046 147454
rect 292810 146898 293046 147134
rect 323530 147218 323766 147454
rect 323530 146898 323766 147134
rect 354250 147218 354486 147454
rect 354250 146898 354486 147134
rect 384970 147218 385206 147454
rect 384970 146898 385206 147134
rect 415690 147218 415926 147454
rect 415690 146898 415926 147134
rect 446410 147218 446646 147454
rect 446410 146898 446646 147134
rect 477130 147218 477366 147454
rect 477130 146898 477366 147134
rect 507850 147218 508086 147454
rect 507850 146898 508086 147134
rect 538570 147218 538806 147454
rect 538570 146898 538806 147134
rect 62410 129218 62646 129454
rect 62410 128898 62646 129134
rect 93130 129218 93366 129454
rect 93130 128898 93366 129134
rect 123850 129218 124086 129454
rect 123850 128898 124086 129134
rect 154570 129218 154806 129454
rect 154570 128898 154806 129134
rect 185290 129218 185526 129454
rect 185290 128898 185526 129134
rect 216010 129218 216246 129454
rect 216010 128898 216246 129134
rect 246730 129218 246966 129454
rect 246730 128898 246966 129134
rect 277450 129218 277686 129454
rect 277450 128898 277686 129134
rect 308170 129218 308406 129454
rect 308170 128898 308406 129134
rect 338890 129218 339126 129454
rect 338890 128898 339126 129134
rect 369610 129218 369846 129454
rect 369610 128898 369846 129134
rect 400330 129218 400566 129454
rect 400330 128898 400566 129134
rect 431050 129218 431286 129454
rect 431050 128898 431286 129134
rect 461770 129218 462006 129454
rect 461770 128898 462006 129134
rect 492490 129218 492726 129454
rect 492490 128898 492726 129134
rect 523210 129218 523446 129454
rect 523210 128898 523446 129134
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 47050 111218 47286 111454
rect 47050 110898 47286 111134
rect 77770 111218 78006 111454
rect 77770 110898 78006 111134
rect 108490 111218 108726 111454
rect 108490 110898 108726 111134
rect 139210 111218 139446 111454
rect 139210 110898 139446 111134
rect 169930 111218 170166 111454
rect 169930 110898 170166 111134
rect 200650 111218 200886 111454
rect 200650 110898 200886 111134
rect 231370 111218 231606 111454
rect 231370 110898 231606 111134
rect 262090 111218 262326 111454
rect 262090 110898 262326 111134
rect 292810 111218 293046 111454
rect 292810 110898 293046 111134
rect 323530 111218 323766 111454
rect 323530 110898 323766 111134
rect 354250 111218 354486 111454
rect 354250 110898 354486 111134
rect 384970 111218 385206 111454
rect 384970 110898 385206 111134
rect 415690 111218 415926 111454
rect 415690 110898 415926 111134
rect 446410 111218 446646 111454
rect 446410 110898 446646 111134
rect 477130 111218 477366 111454
rect 477130 110898 477366 111134
rect 507850 111218 508086 111454
rect 507850 110898 508086 111134
rect 538570 111218 538806 111454
rect 538570 110898 538806 111134
rect 62410 93218 62646 93454
rect 62410 92898 62646 93134
rect 93130 93218 93366 93454
rect 93130 92898 93366 93134
rect 123850 93218 124086 93454
rect 123850 92898 124086 93134
rect 154570 93218 154806 93454
rect 154570 92898 154806 93134
rect 185290 93218 185526 93454
rect 185290 92898 185526 93134
rect 216010 93218 216246 93454
rect 216010 92898 216246 93134
rect 246730 93218 246966 93454
rect 246730 92898 246966 93134
rect 277450 93218 277686 93454
rect 277450 92898 277686 93134
rect 308170 93218 308406 93454
rect 308170 92898 308406 93134
rect 338890 93218 339126 93454
rect 338890 92898 339126 93134
rect 369610 93218 369846 93454
rect 369610 92898 369846 93134
rect 400330 93218 400566 93454
rect 400330 92898 400566 93134
rect 431050 93218 431286 93454
rect 431050 92898 431286 93134
rect 461770 93218 462006 93454
rect 461770 92898 462006 93134
rect 492490 93218 492726 93454
rect 492490 92898 492726 93134
rect 523210 93218 523446 93454
rect 523210 92898 523446 93134
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 47050 75218 47286 75454
rect 47050 74898 47286 75134
rect 77770 75218 78006 75454
rect 77770 74898 78006 75134
rect 108490 75218 108726 75454
rect 108490 74898 108726 75134
rect 139210 75218 139446 75454
rect 139210 74898 139446 75134
rect 169930 75218 170166 75454
rect 169930 74898 170166 75134
rect 200650 75218 200886 75454
rect 200650 74898 200886 75134
rect 231370 75218 231606 75454
rect 231370 74898 231606 75134
rect 262090 75218 262326 75454
rect 262090 74898 262326 75134
rect 292810 75218 293046 75454
rect 292810 74898 293046 75134
rect 323530 75218 323766 75454
rect 323530 74898 323766 75134
rect 354250 75218 354486 75454
rect 354250 74898 354486 75134
rect 384970 75218 385206 75454
rect 384970 74898 385206 75134
rect 415690 75218 415926 75454
rect 415690 74898 415926 75134
rect 446410 75218 446646 75454
rect 446410 74898 446646 75134
rect 477130 75218 477366 75454
rect 477130 74898 477366 75134
rect 507850 75218 508086 75454
rect 507850 74898 508086 75134
rect 538570 75218 538806 75454
rect 538570 74898 538806 75134
rect 62410 57218 62646 57454
rect 62410 56898 62646 57134
rect 93130 57218 93366 57454
rect 93130 56898 93366 57134
rect 123850 57218 124086 57454
rect 123850 56898 124086 57134
rect 154570 57218 154806 57454
rect 154570 56898 154806 57134
rect 185290 57218 185526 57454
rect 185290 56898 185526 57134
rect 216010 57218 216246 57454
rect 216010 56898 216246 57134
rect 246730 57218 246966 57454
rect 246730 56898 246966 57134
rect 277450 57218 277686 57454
rect 277450 56898 277686 57134
rect 308170 57218 308406 57454
rect 308170 56898 308406 57134
rect 338890 57218 339126 57454
rect 338890 56898 339126 57134
rect 369610 57218 369846 57454
rect 369610 56898 369846 57134
rect 400330 57218 400566 57454
rect 400330 56898 400566 57134
rect 431050 57218 431286 57454
rect 431050 56898 431286 57134
rect 461770 57218 462006 57454
rect 461770 56898 462006 57134
rect 492490 57218 492726 57454
rect 492490 56898 492726 57134
rect 523210 57218 523446 57454
rect 523210 56898 523446 57134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 47050 651454
rect 47286 651218 77770 651454
rect 78006 651218 108490 651454
rect 108726 651218 139210 651454
rect 139446 651218 169930 651454
rect 170166 651218 200650 651454
rect 200886 651218 231370 651454
rect 231606 651218 262090 651454
rect 262326 651218 292810 651454
rect 293046 651218 323530 651454
rect 323766 651218 354250 651454
rect 354486 651218 384970 651454
rect 385206 651218 415690 651454
rect 415926 651218 446410 651454
rect 446646 651218 477130 651454
rect 477366 651218 507850 651454
rect 508086 651218 538570 651454
rect 538806 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 47050 651134
rect 47286 650898 77770 651134
rect 78006 650898 108490 651134
rect 108726 650898 139210 651134
rect 139446 650898 169930 651134
rect 170166 650898 200650 651134
rect 200886 650898 231370 651134
rect 231606 650898 262090 651134
rect 262326 650898 292810 651134
rect 293046 650898 323530 651134
rect 323766 650898 354250 651134
rect 354486 650898 384970 651134
rect 385206 650898 415690 651134
rect 415926 650898 446410 651134
rect 446646 650898 477130 651134
rect 477366 650898 507850 651134
rect 508086 650898 538570 651134
rect 538806 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 62410 633454
rect 62646 633218 93130 633454
rect 93366 633218 123850 633454
rect 124086 633218 154570 633454
rect 154806 633218 185290 633454
rect 185526 633218 216010 633454
rect 216246 633218 246730 633454
rect 246966 633218 277450 633454
rect 277686 633218 308170 633454
rect 308406 633218 338890 633454
rect 339126 633218 369610 633454
rect 369846 633218 400330 633454
rect 400566 633218 431050 633454
rect 431286 633218 461770 633454
rect 462006 633218 492490 633454
rect 492726 633218 523210 633454
rect 523446 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 62410 633134
rect 62646 632898 93130 633134
rect 93366 632898 123850 633134
rect 124086 632898 154570 633134
rect 154806 632898 185290 633134
rect 185526 632898 216010 633134
rect 216246 632898 246730 633134
rect 246966 632898 277450 633134
rect 277686 632898 308170 633134
rect 308406 632898 338890 633134
rect 339126 632898 369610 633134
rect 369846 632898 400330 633134
rect 400566 632898 431050 633134
rect 431286 632898 461770 633134
rect 462006 632898 492490 633134
rect 492726 632898 523210 633134
rect 523446 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 47050 615454
rect 47286 615218 77770 615454
rect 78006 615218 108490 615454
rect 108726 615218 139210 615454
rect 139446 615218 169930 615454
rect 170166 615218 200650 615454
rect 200886 615218 231370 615454
rect 231606 615218 262090 615454
rect 262326 615218 292810 615454
rect 293046 615218 323530 615454
rect 323766 615218 354250 615454
rect 354486 615218 384970 615454
rect 385206 615218 415690 615454
rect 415926 615218 446410 615454
rect 446646 615218 477130 615454
rect 477366 615218 507850 615454
rect 508086 615218 538570 615454
rect 538806 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 47050 615134
rect 47286 614898 77770 615134
rect 78006 614898 108490 615134
rect 108726 614898 139210 615134
rect 139446 614898 169930 615134
rect 170166 614898 200650 615134
rect 200886 614898 231370 615134
rect 231606 614898 262090 615134
rect 262326 614898 292810 615134
rect 293046 614898 323530 615134
rect 323766 614898 354250 615134
rect 354486 614898 384970 615134
rect 385206 614898 415690 615134
rect 415926 614898 446410 615134
rect 446646 614898 477130 615134
rect 477366 614898 507850 615134
rect 508086 614898 538570 615134
rect 538806 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 62410 597454
rect 62646 597218 93130 597454
rect 93366 597218 123850 597454
rect 124086 597218 154570 597454
rect 154806 597218 185290 597454
rect 185526 597218 216010 597454
rect 216246 597218 246730 597454
rect 246966 597218 277450 597454
rect 277686 597218 308170 597454
rect 308406 597218 338890 597454
rect 339126 597218 369610 597454
rect 369846 597218 400330 597454
rect 400566 597218 431050 597454
rect 431286 597218 461770 597454
rect 462006 597218 492490 597454
rect 492726 597218 523210 597454
rect 523446 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 62410 597134
rect 62646 596898 93130 597134
rect 93366 596898 123850 597134
rect 124086 596898 154570 597134
rect 154806 596898 185290 597134
rect 185526 596898 216010 597134
rect 216246 596898 246730 597134
rect 246966 596898 277450 597134
rect 277686 596898 308170 597134
rect 308406 596898 338890 597134
rect 339126 596898 369610 597134
rect 369846 596898 400330 597134
rect 400566 596898 431050 597134
rect 431286 596898 461770 597134
rect 462006 596898 492490 597134
rect 492726 596898 523210 597134
rect 523446 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 47050 579454
rect 47286 579218 77770 579454
rect 78006 579218 108490 579454
rect 108726 579218 139210 579454
rect 139446 579218 169930 579454
rect 170166 579218 200650 579454
rect 200886 579218 231370 579454
rect 231606 579218 262090 579454
rect 262326 579218 292810 579454
rect 293046 579218 323530 579454
rect 323766 579218 354250 579454
rect 354486 579218 384970 579454
rect 385206 579218 415690 579454
rect 415926 579218 446410 579454
rect 446646 579218 477130 579454
rect 477366 579218 507850 579454
rect 508086 579218 538570 579454
rect 538806 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 47050 579134
rect 47286 578898 77770 579134
rect 78006 578898 108490 579134
rect 108726 578898 139210 579134
rect 139446 578898 169930 579134
rect 170166 578898 200650 579134
rect 200886 578898 231370 579134
rect 231606 578898 262090 579134
rect 262326 578898 292810 579134
rect 293046 578898 323530 579134
rect 323766 578898 354250 579134
rect 354486 578898 384970 579134
rect 385206 578898 415690 579134
rect 415926 578898 446410 579134
rect 446646 578898 477130 579134
rect 477366 578898 507850 579134
rect 508086 578898 538570 579134
rect 538806 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 62410 561454
rect 62646 561218 93130 561454
rect 93366 561218 123850 561454
rect 124086 561218 154570 561454
rect 154806 561218 185290 561454
rect 185526 561218 216010 561454
rect 216246 561218 246730 561454
rect 246966 561218 277450 561454
rect 277686 561218 308170 561454
rect 308406 561218 338890 561454
rect 339126 561218 369610 561454
rect 369846 561218 400330 561454
rect 400566 561218 431050 561454
rect 431286 561218 461770 561454
rect 462006 561218 492490 561454
rect 492726 561218 523210 561454
rect 523446 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 62410 561134
rect 62646 560898 93130 561134
rect 93366 560898 123850 561134
rect 124086 560898 154570 561134
rect 154806 560898 185290 561134
rect 185526 560898 216010 561134
rect 216246 560898 246730 561134
rect 246966 560898 277450 561134
rect 277686 560898 308170 561134
rect 308406 560898 338890 561134
rect 339126 560898 369610 561134
rect 369846 560898 400330 561134
rect 400566 560898 431050 561134
rect 431286 560898 461770 561134
rect 462006 560898 492490 561134
rect 492726 560898 523210 561134
rect 523446 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 47050 543454
rect 47286 543218 77770 543454
rect 78006 543218 108490 543454
rect 108726 543218 139210 543454
rect 139446 543218 169930 543454
rect 170166 543218 200650 543454
rect 200886 543218 231370 543454
rect 231606 543218 262090 543454
rect 262326 543218 292810 543454
rect 293046 543218 323530 543454
rect 323766 543218 354250 543454
rect 354486 543218 384970 543454
rect 385206 543218 415690 543454
rect 415926 543218 446410 543454
rect 446646 543218 477130 543454
rect 477366 543218 507850 543454
rect 508086 543218 538570 543454
rect 538806 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 47050 543134
rect 47286 542898 77770 543134
rect 78006 542898 108490 543134
rect 108726 542898 139210 543134
rect 139446 542898 169930 543134
rect 170166 542898 200650 543134
rect 200886 542898 231370 543134
rect 231606 542898 262090 543134
rect 262326 542898 292810 543134
rect 293046 542898 323530 543134
rect 323766 542898 354250 543134
rect 354486 542898 384970 543134
rect 385206 542898 415690 543134
rect 415926 542898 446410 543134
rect 446646 542898 477130 543134
rect 477366 542898 507850 543134
rect 508086 542898 538570 543134
rect 538806 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 62410 525454
rect 62646 525218 93130 525454
rect 93366 525218 123850 525454
rect 124086 525218 154570 525454
rect 154806 525218 185290 525454
rect 185526 525218 216010 525454
rect 216246 525218 246730 525454
rect 246966 525218 277450 525454
rect 277686 525218 308170 525454
rect 308406 525218 338890 525454
rect 339126 525218 369610 525454
rect 369846 525218 400330 525454
rect 400566 525218 431050 525454
rect 431286 525218 461770 525454
rect 462006 525218 492490 525454
rect 492726 525218 523210 525454
rect 523446 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 62410 525134
rect 62646 524898 93130 525134
rect 93366 524898 123850 525134
rect 124086 524898 154570 525134
rect 154806 524898 185290 525134
rect 185526 524898 216010 525134
rect 216246 524898 246730 525134
rect 246966 524898 277450 525134
rect 277686 524898 308170 525134
rect 308406 524898 338890 525134
rect 339126 524898 369610 525134
rect 369846 524898 400330 525134
rect 400566 524898 431050 525134
rect 431286 524898 461770 525134
rect 462006 524898 492490 525134
rect 492726 524898 523210 525134
rect 523446 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 47050 507454
rect 47286 507218 77770 507454
rect 78006 507218 108490 507454
rect 108726 507218 139210 507454
rect 139446 507218 169930 507454
rect 170166 507218 200650 507454
rect 200886 507218 231370 507454
rect 231606 507218 262090 507454
rect 262326 507218 292810 507454
rect 293046 507218 323530 507454
rect 323766 507218 354250 507454
rect 354486 507218 384970 507454
rect 385206 507218 415690 507454
rect 415926 507218 446410 507454
rect 446646 507218 477130 507454
rect 477366 507218 507850 507454
rect 508086 507218 538570 507454
rect 538806 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 47050 507134
rect 47286 506898 77770 507134
rect 78006 506898 108490 507134
rect 108726 506898 139210 507134
rect 139446 506898 169930 507134
rect 170166 506898 200650 507134
rect 200886 506898 231370 507134
rect 231606 506898 262090 507134
rect 262326 506898 292810 507134
rect 293046 506898 323530 507134
rect 323766 506898 354250 507134
rect 354486 506898 384970 507134
rect 385206 506898 415690 507134
rect 415926 506898 446410 507134
rect 446646 506898 477130 507134
rect 477366 506898 507850 507134
rect 508086 506898 538570 507134
rect 538806 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 62410 489454
rect 62646 489218 93130 489454
rect 93366 489218 123850 489454
rect 124086 489218 154570 489454
rect 154806 489218 185290 489454
rect 185526 489218 216010 489454
rect 216246 489218 246730 489454
rect 246966 489218 277450 489454
rect 277686 489218 308170 489454
rect 308406 489218 338890 489454
rect 339126 489218 369610 489454
rect 369846 489218 400330 489454
rect 400566 489218 431050 489454
rect 431286 489218 461770 489454
rect 462006 489218 492490 489454
rect 492726 489218 523210 489454
rect 523446 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 62410 489134
rect 62646 488898 93130 489134
rect 93366 488898 123850 489134
rect 124086 488898 154570 489134
rect 154806 488898 185290 489134
rect 185526 488898 216010 489134
rect 216246 488898 246730 489134
rect 246966 488898 277450 489134
rect 277686 488898 308170 489134
rect 308406 488898 338890 489134
rect 339126 488898 369610 489134
rect 369846 488898 400330 489134
rect 400566 488898 431050 489134
rect 431286 488898 461770 489134
rect 462006 488898 492490 489134
rect 492726 488898 523210 489134
rect 523446 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 47050 471454
rect 47286 471218 77770 471454
rect 78006 471218 108490 471454
rect 108726 471218 139210 471454
rect 139446 471218 169930 471454
rect 170166 471218 200650 471454
rect 200886 471218 231370 471454
rect 231606 471218 262090 471454
rect 262326 471218 292810 471454
rect 293046 471218 323530 471454
rect 323766 471218 354250 471454
rect 354486 471218 384970 471454
rect 385206 471218 415690 471454
rect 415926 471218 446410 471454
rect 446646 471218 477130 471454
rect 477366 471218 507850 471454
rect 508086 471218 538570 471454
rect 538806 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 47050 471134
rect 47286 470898 77770 471134
rect 78006 470898 108490 471134
rect 108726 470898 139210 471134
rect 139446 470898 169930 471134
rect 170166 470898 200650 471134
rect 200886 470898 231370 471134
rect 231606 470898 262090 471134
rect 262326 470898 292810 471134
rect 293046 470898 323530 471134
rect 323766 470898 354250 471134
rect 354486 470898 384970 471134
rect 385206 470898 415690 471134
rect 415926 470898 446410 471134
rect 446646 470898 477130 471134
rect 477366 470898 507850 471134
rect 508086 470898 538570 471134
rect 538806 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 62410 453454
rect 62646 453218 93130 453454
rect 93366 453218 123850 453454
rect 124086 453218 154570 453454
rect 154806 453218 185290 453454
rect 185526 453218 216010 453454
rect 216246 453218 246730 453454
rect 246966 453218 277450 453454
rect 277686 453218 308170 453454
rect 308406 453218 338890 453454
rect 339126 453218 369610 453454
rect 369846 453218 400330 453454
rect 400566 453218 431050 453454
rect 431286 453218 461770 453454
rect 462006 453218 492490 453454
rect 492726 453218 523210 453454
rect 523446 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 62410 453134
rect 62646 452898 93130 453134
rect 93366 452898 123850 453134
rect 124086 452898 154570 453134
rect 154806 452898 185290 453134
rect 185526 452898 216010 453134
rect 216246 452898 246730 453134
rect 246966 452898 277450 453134
rect 277686 452898 308170 453134
rect 308406 452898 338890 453134
rect 339126 452898 369610 453134
rect 369846 452898 400330 453134
rect 400566 452898 431050 453134
rect 431286 452898 461770 453134
rect 462006 452898 492490 453134
rect 492726 452898 523210 453134
rect 523446 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 47050 435454
rect 47286 435218 77770 435454
rect 78006 435218 108490 435454
rect 108726 435218 139210 435454
rect 139446 435218 169930 435454
rect 170166 435218 200650 435454
rect 200886 435218 231370 435454
rect 231606 435218 262090 435454
rect 262326 435218 292810 435454
rect 293046 435218 323530 435454
rect 323766 435218 354250 435454
rect 354486 435218 384970 435454
rect 385206 435218 415690 435454
rect 415926 435218 446410 435454
rect 446646 435218 477130 435454
rect 477366 435218 507850 435454
rect 508086 435218 538570 435454
rect 538806 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 47050 435134
rect 47286 434898 77770 435134
rect 78006 434898 108490 435134
rect 108726 434898 139210 435134
rect 139446 434898 169930 435134
rect 170166 434898 200650 435134
rect 200886 434898 231370 435134
rect 231606 434898 262090 435134
rect 262326 434898 292810 435134
rect 293046 434898 323530 435134
rect 323766 434898 354250 435134
rect 354486 434898 384970 435134
rect 385206 434898 415690 435134
rect 415926 434898 446410 435134
rect 446646 434898 477130 435134
rect 477366 434898 507850 435134
rect 508086 434898 538570 435134
rect 538806 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 62410 417454
rect 62646 417218 93130 417454
rect 93366 417218 123850 417454
rect 124086 417218 154570 417454
rect 154806 417218 185290 417454
rect 185526 417218 216010 417454
rect 216246 417218 246730 417454
rect 246966 417218 277450 417454
rect 277686 417218 308170 417454
rect 308406 417218 338890 417454
rect 339126 417218 369610 417454
rect 369846 417218 400330 417454
rect 400566 417218 431050 417454
rect 431286 417218 461770 417454
rect 462006 417218 492490 417454
rect 492726 417218 523210 417454
rect 523446 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 62410 417134
rect 62646 416898 93130 417134
rect 93366 416898 123850 417134
rect 124086 416898 154570 417134
rect 154806 416898 185290 417134
rect 185526 416898 216010 417134
rect 216246 416898 246730 417134
rect 246966 416898 277450 417134
rect 277686 416898 308170 417134
rect 308406 416898 338890 417134
rect 339126 416898 369610 417134
rect 369846 416898 400330 417134
rect 400566 416898 431050 417134
rect 431286 416898 461770 417134
rect 462006 416898 492490 417134
rect 492726 416898 523210 417134
rect 523446 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 47050 399454
rect 47286 399218 77770 399454
rect 78006 399218 108490 399454
rect 108726 399218 139210 399454
rect 139446 399218 169930 399454
rect 170166 399218 200650 399454
rect 200886 399218 231370 399454
rect 231606 399218 262090 399454
rect 262326 399218 292810 399454
rect 293046 399218 323530 399454
rect 323766 399218 354250 399454
rect 354486 399218 384970 399454
rect 385206 399218 415690 399454
rect 415926 399218 446410 399454
rect 446646 399218 477130 399454
rect 477366 399218 507850 399454
rect 508086 399218 538570 399454
rect 538806 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 47050 399134
rect 47286 398898 77770 399134
rect 78006 398898 108490 399134
rect 108726 398898 139210 399134
rect 139446 398898 169930 399134
rect 170166 398898 200650 399134
rect 200886 398898 231370 399134
rect 231606 398898 262090 399134
rect 262326 398898 292810 399134
rect 293046 398898 323530 399134
rect 323766 398898 354250 399134
rect 354486 398898 384970 399134
rect 385206 398898 415690 399134
rect 415926 398898 446410 399134
rect 446646 398898 477130 399134
rect 477366 398898 507850 399134
rect 508086 398898 538570 399134
rect 538806 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 62410 381454
rect 62646 381218 93130 381454
rect 93366 381218 123850 381454
rect 124086 381218 154570 381454
rect 154806 381218 185290 381454
rect 185526 381218 216010 381454
rect 216246 381218 246730 381454
rect 246966 381218 277450 381454
rect 277686 381218 308170 381454
rect 308406 381218 338890 381454
rect 339126 381218 369610 381454
rect 369846 381218 400330 381454
rect 400566 381218 431050 381454
rect 431286 381218 461770 381454
rect 462006 381218 492490 381454
rect 492726 381218 523210 381454
rect 523446 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 62410 381134
rect 62646 380898 93130 381134
rect 93366 380898 123850 381134
rect 124086 380898 154570 381134
rect 154806 380898 185290 381134
rect 185526 380898 216010 381134
rect 216246 380898 246730 381134
rect 246966 380898 277450 381134
rect 277686 380898 308170 381134
rect 308406 380898 338890 381134
rect 339126 380898 369610 381134
rect 369846 380898 400330 381134
rect 400566 380898 431050 381134
rect 431286 380898 461770 381134
rect 462006 380898 492490 381134
rect 492726 380898 523210 381134
rect 523446 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 47050 363454
rect 47286 363218 77770 363454
rect 78006 363218 108490 363454
rect 108726 363218 139210 363454
rect 139446 363218 169930 363454
rect 170166 363218 200650 363454
rect 200886 363218 231370 363454
rect 231606 363218 262090 363454
rect 262326 363218 292810 363454
rect 293046 363218 323530 363454
rect 323766 363218 354250 363454
rect 354486 363218 384970 363454
rect 385206 363218 415690 363454
rect 415926 363218 446410 363454
rect 446646 363218 477130 363454
rect 477366 363218 507850 363454
rect 508086 363218 538570 363454
rect 538806 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 47050 363134
rect 47286 362898 77770 363134
rect 78006 362898 108490 363134
rect 108726 362898 139210 363134
rect 139446 362898 169930 363134
rect 170166 362898 200650 363134
rect 200886 362898 231370 363134
rect 231606 362898 262090 363134
rect 262326 362898 292810 363134
rect 293046 362898 323530 363134
rect 323766 362898 354250 363134
rect 354486 362898 384970 363134
rect 385206 362898 415690 363134
rect 415926 362898 446410 363134
rect 446646 362898 477130 363134
rect 477366 362898 507850 363134
rect 508086 362898 538570 363134
rect 538806 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 62410 345454
rect 62646 345218 93130 345454
rect 93366 345218 123850 345454
rect 124086 345218 154570 345454
rect 154806 345218 185290 345454
rect 185526 345218 216010 345454
rect 216246 345218 246730 345454
rect 246966 345218 277450 345454
rect 277686 345218 308170 345454
rect 308406 345218 338890 345454
rect 339126 345218 369610 345454
rect 369846 345218 400330 345454
rect 400566 345218 431050 345454
rect 431286 345218 461770 345454
rect 462006 345218 492490 345454
rect 492726 345218 523210 345454
rect 523446 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 62410 345134
rect 62646 344898 93130 345134
rect 93366 344898 123850 345134
rect 124086 344898 154570 345134
rect 154806 344898 185290 345134
rect 185526 344898 216010 345134
rect 216246 344898 246730 345134
rect 246966 344898 277450 345134
rect 277686 344898 308170 345134
rect 308406 344898 338890 345134
rect 339126 344898 369610 345134
rect 369846 344898 400330 345134
rect 400566 344898 431050 345134
rect 431286 344898 461770 345134
rect 462006 344898 492490 345134
rect 492726 344898 523210 345134
rect 523446 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 47050 327454
rect 47286 327218 77770 327454
rect 78006 327218 108490 327454
rect 108726 327218 139210 327454
rect 139446 327218 169930 327454
rect 170166 327218 200650 327454
rect 200886 327218 231370 327454
rect 231606 327218 262090 327454
rect 262326 327218 292810 327454
rect 293046 327218 323530 327454
rect 323766 327218 354250 327454
rect 354486 327218 384970 327454
rect 385206 327218 415690 327454
rect 415926 327218 446410 327454
rect 446646 327218 477130 327454
rect 477366 327218 507850 327454
rect 508086 327218 538570 327454
rect 538806 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 47050 327134
rect 47286 326898 77770 327134
rect 78006 326898 108490 327134
rect 108726 326898 139210 327134
rect 139446 326898 169930 327134
rect 170166 326898 200650 327134
rect 200886 326898 231370 327134
rect 231606 326898 262090 327134
rect 262326 326898 292810 327134
rect 293046 326898 323530 327134
rect 323766 326898 354250 327134
rect 354486 326898 384970 327134
rect 385206 326898 415690 327134
rect 415926 326898 446410 327134
rect 446646 326898 477130 327134
rect 477366 326898 507850 327134
rect 508086 326898 538570 327134
rect 538806 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 62410 309454
rect 62646 309218 93130 309454
rect 93366 309218 123850 309454
rect 124086 309218 154570 309454
rect 154806 309218 185290 309454
rect 185526 309218 216010 309454
rect 216246 309218 246730 309454
rect 246966 309218 277450 309454
rect 277686 309218 308170 309454
rect 308406 309218 338890 309454
rect 339126 309218 369610 309454
rect 369846 309218 400330 309454
rect 400566 309218 431050 309454
rect 431286 309218 461770 309454
rect 462006 309218 492490 309454
rect 492726 309218 523210 309454
rect 523446 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 62410 309134
rect 62646 308898 93130 309134
rect 93366 308898 123850 309134
rect 124086 308898 154570 309134
rect 154806 308898 185290 309134
rect 185526 308898 216010 309134
rect 216246 308898 246730 309134
rect 246966 308898 277450 309134
rect 277686 308898 308170 309134
rect 308406 308898 338890 309134
rect 339126 308898 369610 309134
rect 369846 308898 400330 309134
rect 400566 308898 431050 309134
rect 431286 308898 461770 309134
rect 462006 308898 492490 309134
rect 492726 308898 523210 309134
rect 523446 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 47050 291454
rect 47286 291218 77770 291454
rect 78006 291218 108490 291454
rect 108726 291218 139210 291454
rect 139446 291218 169930 291454
rect 170166 291218 200650 291454
rect 200886 291218 231370 291454
rect 231606 291218 262090 291454
rect 262326 291218 292810 291454
rect 293046 291218 323530 291454
rect 323766 291218 354250 291454
rect 354486 291218 384970 291454
rect 385206 291218 415690 291454
rect 415926 291218 446410 291454
rect 446646 291218 477130 291454
rect 477366 291218 507850 291454
rect 508086 291218 538570 291454
rect 538806 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 47050 291134
rect 47286 290898 77770 291134
rect 78006 290898 108490 291134
rect 108726 290898 139210 291134
rect 139446 290898 169930 291134
rect 170166 290898 200650 291134
rect 200886 290898 231370 291134
rect 231606 290898 262090 291134
rect 262326 290898 292810 291134
rect 293046 290898 323530 291134
rect 323766 290898 354250 291134
rect 354486 290898 384970 291134
rect 385206 290898 415690 291134
rect 415926 290898 446410 291134
rect 446646 290898 477130 291134
rect 477366 290898 507850 291134
rect 508086 290898 538570 291134
rect 538806 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 62410 273454
rect 62646 273218 93130 273454
rect 93366 273218 123850 273454
rect 124086 273218 154570 273454
rect 154806 273218 185290 273454
rect 185526 273218 216010 273454
rect 216246 273218 246730 273454
rect 246966 273218 277450 273454
rect 277686 273218 308170 273454
rect 308406 273218 338890 273454
rect 339126 273218 369610 273454
rect 369846 273218 400330 273454
rect 400566 273218 431050 273454
rect 431286 273218 461770 273454
rect 462006 273218 492490 273454
rect 492726 273218 523210 273454
rect 523446 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 62410 273134
rect 62646 272898 93130 273134
rect 93366 272898 123850 273134
rect 124086 272898 154570 273134
rect 154806 272898 185290 273134
rect 185526 272898 216010 273134
rect 216246 272898 246730 273134
rect 246966 272898 277450 273134
rect 277686 272898 308170 273134
rect 308406 272898 338890 273134
rect 339126 272898 369610 273134
rect 369846 272898 400330 273134
rect 400566 272898 431050 273134
rect 431286 272898 461770 273134
rect 462006 272898 492490 273134
rect 492726 272898 523210 273134
rect 523446 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 47050 255454
rect 47286 255218 77770 255454
rect 78006 255218 108490 255454
rect 108726 255218 139210 255454
rect 139446 255218 169930 255454
rect 170166 255218 200650 255454
rect 200886 255218 231370 255454
rect 231606 255218 262090 255454
rect 262326 255218 292810 255454
rect 293046 255218 323530 255454
rect 323766 255218 354250 255454
rect 354486 255218 384970 255454
rect 385206 255218 415690 255454
rect 415926 255218 446410 255454
rect 446646 255218 477130 255454
rect 477366 255218 507850 255454
rect 508086 255218 538570 255454
rect 538806 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 47050 255134
rect 47286 254898 77770 255134
rect 78006 254898 108490 255134
rect 108726 254898 139210 255134
rect 139446 254898 169930 255134
rect 170166 254898 200650 255134
rect 200886 254898 231370 255134
rect 231606 254898 262090 255134
rect 262326 254898 292810 255134
rect 293046 254898 323530 255134
rect 323766 254898 354250 255134
rect 354486 254898 384970 255134
rect 385206 254898 415690 255134
rect 415926 254898 446410 255134
rect 446646 254898 477130 255134
rect 477366 254898 507850 255134
rect 508086 254898 538570 255134
rect 538806 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 62410 237454
rect 62646 237218 93130 237454
rect 93366 237218 123850 237454
rect 124086 237218 154570 237454
rect 154806 237218 185290 237454
rect 185526 237218 216010 237454
rect 216246 237218 246730 237454
rect 246966 237218 277450 237454
rect 277686 237218 308170 237454
rect 308406 237218 338890 237454
rect 339126 237218 369610 237454
rect 369846 237218 400330 237454
rect 400566 237218 431050 237454
rect 431286 237218 461770 237454
rect 462006 237218 492490 237454
rect 492726 237218 523210 237454
rect 523446 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 62410 237134
rect 62646 236898 93130 237134
rect 93366 236898 123850 237134
rect 124086 236898 154570 237134
rect 154806 236898 185290 237134
rect 185526 236898 216010 237134
rect 216246 236898 246730 237134
rect 246966 236898 277450 237134
rect 277686 236898 308170 237134
rect 308406 236898 338890 237134
rect 339126 236898 369610 237134
rect 369846 236898 400330 237134
rect 400566 236898 431050 237134
rect 431286 236898 461770 237134
rect 462006 236898 492490 237134
rect 492726 236898 523210 237134
rect 523446 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 47050 219454
rect 47286 219218 77770 219454
rect 78006 219218 108490 219454
rect 108726 219218 139210 219454
rect 139446 219218 169930 219454
rect 170166 219218 200650 219454
rect 200886 219218 231370 219454
rect 231606 219218 262090 219454
rect 262326 219218 292810 219454
rect 293046 219218 323530 219454
rect 323766 219218 354250 219454
rect 354486 219218 384970 219454
rect 385206 219218 415690 219454
rect 415926 219218 446410 219454
rect 446646 219218 477130 219454
rect 477366 219218 507850 219454
rect 508086 219218 538570 219454
rect 538806 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 47050 219134
rect 47286 218898 77770 219134
rect 78006 218898 108490 219134
rect 108726 218898 139210 219134
rect 139446 218898 169930 219134
rect 170166 218898 200650 219134
rect 200886 218898 231370 219134
rect 231606 218898 262090 219134
rect 262326 218898 292810 219134
rect 293046 218898 323530 219134
rect 323766 218898 354250 219134
rect 354486 218898 384970 219134
rect 385206 218898 415690 219134
rect 415926 218898 446410 219134
rect 446646 218898 477130 219134
rect 477366 218898 507850 219134
rect 508086 218898 538570 219134
rect 538806 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 62410 201454
rect 62646 201218 93130 201454
rect 93366 201218 123850 201454
rect 124086 201218 154570 201454
rect 154806 201218 185290 201454
rect 185526 201218 216010 201454
rect 216246 201218 246730 201454
rect 246966 201218 277450 201454
rect 277686 201218 308170 201454
rect 308406 201218 338890 201454
rect 339126 201218 369610 201454
rect 369846 201218 400330 201454
rect 400566 201218 431050 201454
rect 431286 201218 461770 201454
rect 462006 201218 492490 201454
rect 492726 201218 523210 201454
rect 523446 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 62410 201134
rect 62646 200898 93130 201134
rect 93366 200898 123850 201134
rect 124086 200898 154570 201134
rect 154806 200898 185290 201134
rect 185526 200898 216010 201134
rect 216246 200898 246730 201134
rect 246966 200898 277450 201134
rect 277686 200898 308170 201134
rect 308406 200898 338890 201134
rect 339126 200898 369610 201134
rect 369846 200898 400330 201134
rect 400566 200898 431050 201134
rect 431286 200898 461770 201134
rect 462006 200898 492490 201134
rect 492726 200898 523210 201134
rect 523446 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 47050 183454
rect 47286 183218 77770 183454
rect 78006 183218 108490 183454
rect 108726 183218 139210 183454
rect 139446 183218 169930 183454
rect 170166 183218 200650 183454
rect 200886 183218 231370 183454
rect 231606 183218 262090 183454
rect 262326 183218 292810 183454
rect 293046 183218 323530 183454
rect 323766 183218 354250 183454
rect 354486 183218 384970 183454
rect 385206 183218 415690 183454
rect 415926 183218 446410 183454
rect 446646 183218 477130 183454
rect 477366 183218 507850 183454
rect 508086 183218 538570 183454
rect 538806 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 47050 183134
rect 47286 182898 77770 183134
rect 78006 182898 108490 183134
rect 108726 182898 139210 183134
rect 139446 182898 169930 183134
rect 170166 182898 200650 183134
rect 200886 182898 231370 183134
rect 231606 182898 262090 183134
rect 262326 182898 292810 183134
rect 293046 182898 323530 183134
rect 323766 182898 354250 183134
rect 354486 182898 384970 183134
rect 385206 182898 415690 183134
rect 415926 182898 446410 183134
rect 446646 182898 477130 183134
rect 477366 182898 507850 183134
rect 508086 182898 538570 183134
rect 538806 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 62410 165454
rect 62646 165218 93130 165454
rect 93366 165218 123850 165454
rect 124086 165218 154570 165454
rect 154806 165218 185290 165454
rect 185526 165218 216010 165454
rect 216246 165218 246730 165454
rect 246966 165218 277450 165454
rect 277686 165218 308170 165454
rect 308406 165218 338890 165454
rect 339126 165218 369610 165454
rect 369846 165218 400330 165454
rect 400566 165218 431050 165454
rect 431286 165218 461770 165454
rect 462006 165218 492490 165454
rect 492726 165218 523210 165454
rect 523446 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 62410 165134
rect 62646 164898 93130 165134
rect 93366 164898 123850 165134
rect 124086 164898 154570 165134
rect 154806 164898 185290 165134
rect 185526 164898 216010 165134
rect 216246 164898 246730 165134
rect 246966 164898 277450 165134
rect 277686 164898 308170 165134
rect 308406 164898 338890 165134
rect 339126 164898 369610 165134
rect 369846 164898 400330 165134
rect 400566 164898 431050 165134
rect 431286 164898 461770 165134
rect 462006 164898 492490 165134
rect 492726 164898 523210 165134
rect 523446 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 47050 147454
rect 47286 147218 77770 147454
rect 78006 147218 108490 147454
rect 108726 147218 139210 147454
rect 139446 147218 169930 147454
rect 170166 147218 200650 147454
rect 200886 147218 231370 147454
rect 231606 147218 262090 147454
rect 262326 147218 292810 147454
rect 293046 147218 323530 147454
rect 323766 147218 354250 147454
rect 354486 147218 384970 147454
rect 385206 147218 415690 147454
rect 415926 147218 446410 147454
rect 446646 147218 477130 147454
rect 477366 147218 507850 147454
rect 508086 147218 538570 147454
rect 538806 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 47050 147134
rect 47286 146898 77770 147134
rect 78006 146898 108490 147134
rect 108726 146898 139210 147134
rect 139446 146898 169930 147134
rect 170166 146898 200650 147134
rect 200886 146898 231370 147134
rect 231606 146898 262090 147134
rect 262326 146898 292810 147134
rect 293046 146898 323530 147134
rect 323766 146898 354250 147134
rect 354486 146898 384970 147134
rect 385206 146898 415690 147134
rect 415926 146898 446410 147134
rect 446646 146898 477130 147134
rect 477366 146898 507850 147134
rect 508086 146898 538570 147134
rect 538806 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 62410 129454
rect 62646 129218 93130 129454
rect 93366 129218 123850 129454
rect 124086 129218 154570 129454
rect 154806 129218 185290 129454
rect 185526 129218 216010 129454
rect 216246 129218 246730 129454
rect 246966 129218 277450 129454
rect 277686 129218 308170 129454
rect 308406 129218 338890 129454
rect 339126 129218 369610 129454
rect 369846 129218 400330 129454
rect 400566 129218 431050 129454
rect 431286 129218 461770 129454
rect 462006 129218 492490 129454
rect 492726 129218 523210 129454
rect 523446 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 62410 129134
rect 62646 128898 93130 129134
rect 93366 128898 123850 129134
rect 124086 128898 154570 129134
rect 154806 128898 185290 129134
rect 185526 128898 216010 129134
rect 216246 128898 246730 129134
rect 246966 128898 277450 129134
rect 277686 128898 308170 129134
rect 308406 128898 338890 129134
rect 339126 128898 369610 129134
rect 369846 128898 400330 129134
rect 400566 128898 431050 129134
rect 431286 128898 461770 129134
rect 462006 128898 492490 129134
rect 492726 128898 523210 129134
rect 523446 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 47050 111454
rect 47286 111218 77770 111454
rect 78006 111218 108490 111454
rect 108726 111218 139210 111454
rect 139446 111218 169930 111454
rect 170166 111218 200650 111454
rect 200886 111218 231370 111454
rect 231606 111218 262090 111454
rect 262326 111218 292810 111454
rect 293046 111218 323530 111454
rect 323766 111218 354250 111454
rect 354486 111218 384970 111454
rect 385206 111218 415690 111454
rect 415926 111218 446410 111454
rect 446646 111218 477130 111454
rect 477366 111218 507850 111454
rect 508086 111218 538570 111454
rect 538806 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 47050 111134
rect 47286 110898 77770 111134
rect 78006 110898 108490 111134
rect 108726 110898 139210 111134
rect 139446 110898 169930 111134
rect 170166 110898 200650 111134
rect 200886 110898 231370 111134
rect 231606 110898 262090 111134
rect 262326 110898 292810 111134
rect 293046 110898 323530 111134
rect 323766 110898 354250 111134
rect 354486 110898 384970 111134
rect 385206 110898 415690 111134
rect 415926 110898 446410 111134
rect 446646 110898 477130 111134
rect 477366 110898 507850 111134
rect 508086 110898 538570 111134
rect 538806 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 62410 93454
rect 62646 93218 93130 93454
rect 93366 93218 123850 93454
rect 124086 93218 154570 93454
rect 154806 93218 185290 93454
rect 185526 93218 216010 93454
rect 216246 93218 246730 93454
rect 246966 93218 277450 93454
rect 277686 93218 308170 93454
rect 308406 93218 338890 93454
rect 339126 93218 369610 93454
rect 369846 93218 400330 93454
rect 400566 93218 431050 93454
rect 431286 93218 461770 93454
rect 462006 93218 492490 93454
rect 492726 93218 523210 93454
rect 523446 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 62410 93134
rect 62646 92898 93130 93134
rect 93366 92898 123850 93134
rect 124086 92898 154570 93134
rect 154806 92898 185290 93134
rect 185526 92898 216010 93134
rect 216246 92898 246730 93134
rect 246966 92898 277450 93134
rect 277686 92898 308170 93134
rect 308406 92898 338890 93134
rect 339126 92898 369610 93134
rect 369846 92898 400330 93134
rect 400566 92898 431050 93134
rect 431286 92898 461770 93134
rect 462006 92898 492490 93134
rect 492726 92898 523210 93134
rect 523446 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 47050 75454
rect 47286 75218 77770 75454
rect 78006 75218 108490 75454
rect 108726 75218 139210 75454
rect 139446 75218 169930 75454
rect 170166 75218 200650 75454
rect 200886 75218 231370 75454
rect 231606 75218 262090 75454
rect 262326 75218 292810 75454
rect 293046 75218 323530 75454
rect 323766 75218 354250 75454
rect 354486 75218 384970 75454
rect 385206 75218 415690 75454
rect 415926 75218 446410 75454
rect 446646 75218 477130 75454
rect 477366 75218 507850 75454
rect 508086 75218 538570 75454
rect 538806 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 47050 75134
rect 47286 74898 77770 75134
rect 78006 74898 108490 75134
rect 108726 74898 139210 75134
rect 139446 74898 169930 75134
rect 170166 74898 200650 75134
rect 200886 74898 231370 75134
rect 231606 74898 262090 75134
rect 262326 74898 292810 75134
rect 293046 74898 323530 75134
rect 323766 74898 354250 75134
rect 354486 74898 384970 75134
rect 385206 74898 415690 75134
rect 415926 74898 446410 75134
rect 446646 74898 477130 75134
rect 477366 74898 507850 75134
rect 508086 74898 538570 75134
rect 538806 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 62410 57454
rect 62646 57218 93130 57454
rect 93366 57218 123850 57454
rect 124086 57218 154570 57454
rect 154806 57218 185290 57454
rect 185526 57218 216010 57454
rect 216246 57218 246730 57454
rect 246966 57218 277450 57454
rect 277686 57218 308170 57454
rect 308406 57218 338890 57454
rect 339126 57218 369610 57454
rect 369846 57218 400330 57454
rect 400566 57218 431050 57454
rect 431286 57218 461770 57454
rect 462006 57218 492490 57454
rect 492726 57218 523210 57454
rect 523446 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 62410 57134
rect 62646 56898 93130 57134
rect 93366 56898 123850 57134
rect 124086 56898 154570 57134
rect 154806 56898 185290 57134
rect 185526 56898 216010 57134
rect 216246 56898 246730 57134
rect 246966 56898 277450 57134
rect 277686 56898 308170 57134
rect 308406 56898 338890 57134
rect 339126 56898 369610 57134
rect 369846 56898 400330 57134
rect 400566 56898 431050 57134
rect 431286 56898 461770 57134
rect 462006 56898 492490 57134
rect 492726 56898 523210 57134
rect 523446 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1641015008
transform 1 0 42800 0 1 53000
box 474 0 500282 602697
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 51000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 657697 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 657697 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 657697 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 657697 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 657697 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 657697 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 657697 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 657697 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 657697 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 657697 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 657697 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 657697 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 657697 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 657697 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 51000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 657697 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 657697 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 657697 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 657697 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 657697 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 657697 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 657697 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 657697 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 657697 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 657697 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 657697 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 657697 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 657697 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 657697 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 657697 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 51000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 657697 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 657697 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 657697 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 657697 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 657697 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 657697 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 657697 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 657697 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 657697 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 657697 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 657697 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 657697 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 657697 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 657697 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 51000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 657697 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 657697 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 657697 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 657697 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 657697 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 657697 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 657697 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 657697 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 657697 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 657697 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 657697 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 657697 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 657697 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 657697 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 51000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 657697 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 657697 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 657697 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 657697 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 657697 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 657697 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 657697 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 657697 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 657697 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 657697 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 657697 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 657697 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 657697 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 657697 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 51000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 657697 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 657697 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 657697 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 657697 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 657697 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 657697 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 657697 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 657697 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 657697 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 657697 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 657697 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 657697 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 657697 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 657697 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 51000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 657697 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 657697 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 657697 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 657697 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 657697 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 657697 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 657697 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 657697 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 657697 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 657697 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 657697 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 657697 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 657697 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 657697 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 51000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 657697 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 657697 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 657697 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 657697 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 657697 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 657697 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 657697 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 657697 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 657697 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 657697 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 657697 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 657697 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 657697 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 657697 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
