magic
tech sky130A
magscale 1 2
timestamp 1641138818
<< obsli1 >>
rect 1104 1445 499991 600049
<< obsm1 >>
rect 474 1436 500282 600080
<< metal2 >>
rect 2134 601897 2190 602697
rect 6458 601897 6514 602697
rect 10874 601897 10930 602697
rect 15290 601897 15346 602697
rect 19706 601897 19762 602697
rect 24030 601897 24086 602697
rect 28446 601897 28502 602697
rect 32862 601897 32918 602697
rect 37278 601897 37334 602697
rect 41602 601897 41658 602697
rect 46018 601897 46074 602697
rect 50434 601897 50490 602697
rect 54850 601897 54906 602697
rect 59174 601897 59230 602697
rect 63590 601897 63646 602697
rect 68006 601897 68062 602697
rect 72422 601897 72478 602697
rect 76746 601897 76802 602697
rect 81162 601897 81218 602697
rect 85578 601897 85634 602697
rect 89994 601897 90050 602697
rect 94318 601897 94374 602697
rect 98734 601897 98790 602697
rect 103150 601897 103206 602697
rect 107566 601897 107622 602697
rect 111890 601897 111946 602697
rect 116306 601897 116362 602697
rect 120722 601897 120778 602697
rect 125138 601897 125194 602697
rect 129462 601897 129518 602697
rect 133878 601897 133934 602697
rect 138294 601897 138350 602697
rect 142710 601897 142766 602697
rect 147034 601897 147090 602697
rect 151450 601897 151506 602697
rect 155866 601897 155922 602697
rect 160282 601897 160338 602697
rect 164606 601897 164662 602697
rect 169022 601897 169078 602697
rect 173438 601897 173494 602697
rect 177854 601897 177910 602697
rect 182178 601897 182234 602697
rect 186594 601897 186650 602697
rect 191010 601897 191066 602697
rect 195426 601897 195482 602697
rect 199750 601897 199806 602697
rect 204166 601897 204222 602697
rect 208582 601897 208638 602697
rect 212998 601897 213054 602697
rect 217322 601897 217378 602697
rect 221738 601897 221794 602697
rect 226154 601897 226210 602697
rect 230570 601897 230626 602697
rect 234894 601897 234950 602697
rect 239310 601897 239366 602697
rect 243726 601897 243782 602697
rect 248142 601897 248198 602697
rect 252558 601897 252614 602697
rect 256882 601897 256938 602697
rect 261298 601897 261354 602697
rect 265714 601897 265770 602697
rect 270130 601897 270186 602697
rect 274454 601897 274510 602697
rect 278870 601897 278926 602697
rect 283286 601897 283342 602697
rect 287702 601897 287758 602697
rect 292026 601897 292082 602697
rect 296442 601897 296498 602697
rect 300858 601897 300914 602697
rect 305274 601897 305330 602697
rect 309598 601897 309654 602697
rect 314014 601897 314070 602697
rect 318430 601897 318486 602697
rect 322846 601897 322902 602697
rect 327170 601897 327226 602697
rect 331586 601897 331642 602697
rect 336002 601897 336058 602697
rect 340418 601897 340474 602697
rect 344742 601897 344798 602697
rect 349158 601897 349214 602697
rect 353574 601897 353630 602697
rect 357990 601897 358046 602697
rect 362314 601897 362370 602697
rect 366730 601897 366786 602697
rect 371146 601897 371202 602697
rect 375562 601897 375618 602697
rect 379886 601897 379942 602697
rect 384302 601897 384358 602697
rect 388718 601897 388774 602697
rect 393134 601897 393190 602697
rect 397458 601897 397514 602697
rect 401874 601897 401930 602697
rect 406290 601897 406346 602697
rect 410706 601897 410762 602697
rect 415030 601897 415086 602697
rect 419446 601897 419502 602697
rect 423862 601897 423918 602697
rect 428278 601897 428334 602697
rect 432602 601897 432658 602697
rect 437018 601897 437074 602697
rect 441434 601897 441490 602697
rect 445850 601897 445906 602697
rect 450174 601897 450230 602697
rect 454590 601897 454646 602697
rect 459006 601897 459062 602697
rect 463422 601897 463478 602697
rect 467746 601897 467802 602697
rect 472162 601897 472218 602697
rect 476578 601897 476634 602697
rect 480994 601897 481050 602697
rect 485318 601897 485374 602697
rect 489734 601897 489790 602697
rect 494150 601897 494206 602697
rect 498566 601897 498622 602697
rect 478 0 534 800
rect 1490 0 1546 800
rect 2502 0 2558 800
rect 3514 0 3570 800
rect 4526 0 4582 800
rect 5538 0 5594 800
rect 6550 0 6606 800
rect 7562 0 7618 800
rect 8574 0 8630 800
rect 9586 0 9642 800
rect 10598 0 10654 800
rect 11610 0 11666 800
rect 12622 0 12678 800
rect 13634 0 13690 800
rect 14646 0 14702 800
rect 15658 0 15714 800
rect 16670 0 16726 800
rect 17682 0 17738 800
rect 18694 0 18750 800
rect 19706 0 19762 800
rect 20718 0 20774 800
rect 21730 0 21786 800
rect 22742 0 22798 800
rect 23754 0 23810 800
rect 24858 0 24914 800
rect 25870 0 25926 800
rect 26882 0 26938 800
rect 27894 0 27950 800
rect 28906 0 28962 800
rect 29918 0 29974 800
rect 30930 0 30986 800
rect 31942 0 31998 800
rect 32954 0 33010 800
rect 33966 0 34022 800
rect 34978 0 35034 800
rect 35990 0 36046 800
rect 37002 0 37058 800
rect 38014 0 38070 800
rect 39026 0 39082 800
rect 40038 0 40094 800
rect 41050 0 41106 800
rect 42062 0 42118 800
rect 43074 0 43130 800
rect 44086 0 44142 800
rect 45098 0 45154 800
rect 46110 0 46166 800
rect 47122 0 47178 800
rect 48226 0 48282 800
rect 49238 0 49294 800
rect 50250 0 50306 800
rect 51262 0 51318 800
rect 52274 0 52330 800
rect 53286 0 53342 800
rect 54298 0 54354 800
rect 55310 0 55366 800
rect 56322 0 56378 800
rect 57334 0 57390 800
rect 58346 0 58402 800
rect 59358 0 59414 800
rect 60370 0 60426 800
rect 61382 0 61438 800
rect 62394 0 62450 800
rect 63406 0 63462 800
rect 64418 0 64474 800
rect 65430 0 65486 800
rect 66442 0 66498 800
rect 67454 0 67510 800
rect 68466 0 68522 800
rect 69478 0 69534 800
rect 70490 0 70546 800
rect 71502 0 71558 800
rect 72606 0 72662 800
rect 73618 0 73674 800
rect 74630 0 74686 800
rect 75642 0 75698 800
rect 76654 0 76710 800
rect 77666 0 77722 800
rect 78678 0 78734 800
rect 79690 0 79746 800
rect 80702 0 80758 800
rect 81714 0 81770 800
rect 82726 0 82782 800
rect 83738 0 83794 800
rect 84750 0 84806 800
rect 85762 0 85818 800
rect 86774 0 86830 800
rect 87786 0 87842 800
rect 88798 0 88854 800
rect 89810 0 89866 800
rect 90822 0 90878 800
rect 91834 0 91890 800
rect 92846 0 92902 800
rect 93858 0 93914 800
rect 94870 0 94926 800
rect 95974 0 96030 800
rect 96986 0 97042 800
rect 97998 0 98054 800
rect 99010 0 99066 800
rect 100022 0 100078 800
rect 101034 0 101090 800
rect 102046 0 102102 800
rect 103058 0 103114 800
rect 104070 0 104126 800
rect 105082 0 105138 800
rect 106094 0 106150 800
rect 107106 0 107162 800
rect 108118 0 108174 800
rect 109130 0 109186 800
rect 110142 0 110198 800
rect 111154 0 111210 800
rect 112166 0 112222 800
rect 113178 0 113234 800
rect 114190 0 114246 800
rect 115202 0 115258 800
rect 116214 0 116270 800
rect 117226 0 117282 800
rect 118238 0 118294 800
rect 119250 0 119306 800
rect 120354 0 120410 800
rect 121366 0 121422 800
rect 122378 0 122434 800
rect 123390 0 123446 800
rect 124402 0 124458 800
rect 125414 0 125470 800
rect 126426 0 126482 800
rect 127438 0 127494 800
rect 128450 0 128506 800
rect 129462 0 129518 800
rect 130474 0 130530 800
rect 131486 0 131542 800
rect 132498 0 132554 800
rect 133510 0 133566 800
rect 134522 0 134578 800
rect 135534 0 135590 800
rect 136546 0 136602 800
rect 137558 0 137614 800
rect 138570 0 138626 800
rect 139582 0 139638 800
rect 140594 0 140650 800
rect 141606 0 141662 800
rect 142618 0 142674 800
rect 143722 0 143778 800
rect 144734 0 144790 800
rect 145746 0 145802 800
rect 146758 0 146814 800
rect 147770 0 147826 800
rect 148782 0 148838 800
rect 149794 0 149850 800
rect 150806 0 150862 800
rect 151818 0 151874 800
rect 152830 0 152886 800
rect 153842 0 153898 800
rect 154854 0 154910 800
rect 155866 0 155922 800
rect 156878 0 156934 800
rect 157890 0 157946 800
rect 158902 0 158958 800
rect 159914 0 159970 800
rect 160926 0 160982 800
rect 161938 0 161994 800
rect 162950 0 163006 800
rect 163962 0 164018 800
rect 164974 0 165030 800
rect 165986 0 166042 800
rect 166998 0 167054 800
rect 168102 0 168158 800
rect 169114 0 169170 800
rect 170126 0 170182 800
rect 171138 0 171194 800
rect 172150 0 172206 800
rect 173162 0 173218 800
rect 174174 0 174230 800
rect 175186 0 175242 800
rect 176198 0 176254 800
rect 177210 0 177266 800
rect 178222 0 178278 800
rect 179234 0 179290 800
rect 180246 0 180302 800
rect 181258 0 181314 800
rect 182270 0 182326 800
rect 183282 0 183338 800
rect 184294 0 184350 800
rect 185306 0 185362 800
rect 186318 0 186374 800
rect 187330 0 187386 800
rect 188342 0 188398 800
rect 189354 0 189410 800
rect 190366 0 190422 800
rect 191470 0 191526 800
rect 192482 0 192538 800
rect 193494 0 193550 800
rect 194506 0 194562 800
rect 195518 0 195574 800
rect 196530 0 196586 800
rect 197542 0 197598 800
rect 198554 0 198610 800
rect 199566 0 199622 800
rect 200578 0 200634 800
rect 201590 0 201646 800
rect 202602 0 202658 800
rect 203614 0 203670 800
rect 204626 0 204682 800
rect 205638 0 205694 800
rect 206650 0 206706 800
rect 207662 0 207718 800
rect 208674 0 208730 800
rect 209686 0 209742 800
rect 210698 0 210754 800
rect 211710 0 211766 800
rect 212722 0 212778 800
rect 213734 0 213790 800
rect 214746 0 214802 800
rect 215850 0 215906 800
rect 216862 0 216918 800
rect 217874 0 217930 800
rect 218886 0 218942 800
rect 219898 0 219954 800
rect 220910 0 220966 800
rect 221922 0 221978 800
rect 222934 0 222990 800
rect 223946 0 224002 800
rect 224958 0 225014 800
rect 225970 0 226026 800
rect 226982 0 227038 800
rect 227994 0 228050 800
rect 229006 0 229062 800
rect 230018 0 230074 800
rect 231030 0 231086 800
rect 232042 0 232098 800
rect 233054 0 233110 800
rect 234066 0 234122 800
rect 235078 0 235134 800
rect 236090 0 236146 800
rect 237102 0 237158 800
rect 238114 0 238170 800
rect 239218 0 239274 800
rect 240230 0 240286 800
rect 241242 0 241298 800
rect 242254 0 242310 800
rect 243266 0 243322 800
rect 244278 0 244334 800
rect 245290 0 245346 800
rect 246302 0 246358 800
rect 247314 0 247370 800
rect 248326 0 248382 800
rect 249338 0 249394 800
rect 250350 0 250406 800
rect 251362 0 251418 800
rect 252374 0 252430 800
rect 253386 0 253442 800
rect 254398 0 254454 800
rect 255410 0 255466 800
rect 256422 0 256478 800
rect 257434 0 257490 800
rect 258446 0 258502 800
rect 259458 0 259514 800
rect 260470 0 260526 800
rect 261482 0 261538 800
rect 262494 0 262550 800
rect 263598 0 263654 800
rect 264610 0 264666 800
rect 265622 0 265678 800
rect 266634 0 266690 800
rect 267646 0 267702 800
rect 268658 0 268714 800
rect 269670 0 269726 800
rect 270682 0 270738 800
rect 271694 0 271750 800
rect 272706 0 272762 800
rect 273718 0 273774 800
rect 274730 0 274786 800
rect 275742 0 275798 800
rect 276754 0 276810 800
rect 277766 0 277822 800
rect 278778 0 278834 800
rect 279790 0 279846 800
rect 280802 0 280858 800
rect 281814 0 281870 800
rect 282826 0 282882 800
rect 283838 0 283894 800
rect 284850 0 284906 800
rect 285862 0 285918 800
rect 286966 0 287022 800
rect 287978 0 288034 800
rect 288990 0 289046 800
rect 290002 0 290058 800
rect 291014 0 291070 800
rect 292026 0 292082 800
rect 293038 0 293094 800
rect 294050 0 294106 800
rect 295062 0 295118 800
rect 296074 0 296130 800
rect 297086 0 297142 800
rect 298098 0 298154 800
rect 299110 0 299166 800
rect 300122 0 300178 800
rect 301134 0 301190 800
rect 302146 0 302202 800
rect 303158 0 303214 800
rect 304170 0 304226 800
rect 305182 0 305238 800
rect 306194 0 306250 800
rect 307206 0 307262 800
rect 308218 0 308274 800
rect 309230 0 309286 800
rect 310242 0 310298 800
rect 311346 0 311402 800
rect 312358 0 312414 800
rect 313370 0 313426 800
rect 314382 0 314438 800
rect 315394 0 315450 800
rect 316406 0 316462 800
rect 317418 0 317474 800
rect 318430 0 318486 800
rect 319442 0 319498 800
rect 320454 0 320510 800
rect 321466 0 321522 800
rect 322478 0 322534 800
rect 323490 0 323546 800
rect 324502 0 324558 800
rect 325514 0 325570 800
rect 326526 0 326582 800
rect 327538 0 327594 800
rect 328550 0 328606 800
rect 329562 0 329618 800
rect 330574 0 330630 800
rect 331586 0 331642 800
rect 332598 0 332654 800
rect 333610 0 333666 800
rect 334714 0 334770 800
rect 335726 0 335782 800
rect 336738 0 336794 800
rect 337750 0 337806 800
rect 338762 0 338818 800
rect 339774 0 339830 800
rect 340786 0 340842 800
rect 341798 0 341854 800
rect 342810 0 342866 800
rect 343822 0 343878 800
rect 344834 0 344890 800
rect 345846 0 345902 800
rect 346858 0 346914 800
rect 347870 0 347926 800
rect 348882 0 348938 800
rect 349894 0 349950 800
rect 350906 0 350962 800
rect 351918 0 351974 800
rect 352930 0 352986 800
rect 353942 0 353998 800
rect 354954 0 355010 800
rect 355966 0 356022 800
rect 356978 0 357034 800
rect 357990 0 358046 800
rect 359094 0 359150 800
rect 360106 0 360162 800
rect 361118 0 361174 800
rect 362130 0 362186 800
rect 363142 0 363198 800
rect 364154 0 364210 800
rect 365166 0 365222 800
rect 366178 0 366234 800
rect 367190 0 367246 800
rect 368202 0 368258 800
rect 369214 0 369270 800
rect 370226 0 370282 800
rect 371238 0 371294 800
rect 372250 0 372306 800
rect 373262 0 373318 800
rect 374274 0 374330 800
rect 375286 0 375342 800
rect 376298 0 376354 800
rect 377310 0 377366 800
rect 378322 0 378378 800
rect 379334 0 379390 800
rect 380346 0 380402 800
rect 381358 0 381414 800
rect 382462 0 382518 800
rect 383474 0 383530 800
rect 384486 0 384542 800
rect 385498 0 385554 800
rect 386510 0 386566 800
rect 387522 0 387578 800
rect 388534 0 388590 800
rect 389546 0 389602 800
rect 390558 0 390614 800
rect 391570 0 391626 800
rect 392582 0 392638 800
rect 393594 0 393650 800
rect 394606 0 394662 800
rect 395618 0 395674 800
rect 396630 0 396686 800
rect 397642 0 397698 800
rect 398654 0 398710 800
rect 399666 0 399722 800
rect 400678 0 400734 800
rect 401690 0 401746 800
rect 402702 0 402758 800
rect 403714 0 403770 800
rect 404726 0 404782 800
rect 405738 0 405794 800
rect 406842 0 406898 800
rect 407854 0 407910 800
rect 408866 0 408922 800
rect 409878 0 409934 800
rect 410890 0 410946 800
rect 411902 0 411958 800
rect 412914 0 412970 800
rect 413926 0 413982 800
rect 414938 0 414994 800
rect 415950 0 416006 800
rect 416962 0 417018 800
rect 417974 0 418030 800
rect 418986 0 419042 800
rect 419998 0 420054 800
rect 421010 0 421066 800
rect 422022 0 422078 800
rect 423034 0 423090 800
rect 424046 0 424102 800
rect 425058 0 425114 800
rect 426070 0 426126 800
rect 427082 0 427138 800
rect 428094 0 428150 800
rect 429106 0 429162 800
rect 430210 0 430266 800
rect 431222 0 431278 800
rect 432234 0 432290 800
rect 433246 0 433302 800
rect 434258 0 434314 800
rect 435270 0 435326 800
rect 436282 0 436338 800
rect 437294 0 437350 800
rect 438306 0 438362 800
rect 439318 0 439374 800
rect 440330 0 440386 800
rect 441342 0 441398 800
rect 442354 0 442410 800
rect 443366 0 443422 800
rect 444378 0 444434 800
rect 445390 0 445446 800
rect 446402 0 446458 800
rect 447414 0 447470 800
rect 448426 0 448482 800
rect 449438 0 449494 800
rect 450450 0 450506 800
rect 451462 0 451518 800
rect 452474 0 452530 800
rect 453486 0 453542 800
rect 454590 0 454646 800
rect 455602 0 455658 800
rect 456614 0 456670 800
rect 457626 0 457682 800
rect 458638 0 458694 800
rect 459650 0 459706 800
rect 460662 0 460718 800
rect 461674 0 461730 800
rect 462686 0 462742 800
rect 463698 0 463754 800
rect 464710 0 464766 800
rect 465722 0 465778 800
rect 466734 0 466790 800
rect 467746 0 467802 800
rect 468758 0 468814 800
rect 469770 0 469826 800
rect 470782 0 470838 800
rect 471794 0 471850 800
rect 472806 0 472862 800
rect 473818 0 473874 800
rect 474830 0 474886 800
rect 475842 0 475898 800
rect 476854 0 476910 800
rect 477958 0 478014 800
rect 478970 0 479026 800
rect 479982 0 480038 800
rect 480994 0 481050 800
rect 482006 0 482062 800
rect 483018 0 483074 800
rect 484030 0 484086 800
rect 485042 0 485098 800
rect 486054 0 486110 800
rect 487066 0 487122 800
rect 488078 0 488134 800
rect 489090 0 489146 800
rect 490102 0 490158 800
rect 491114 0 491170 800
rect 492126 0 492182 800
rect 493138 0 493194 800
rect 494150 0 494206 800
rect 495162 0 495218 800
rect 496174 0 496230 800
rect 497186 0 497242 800
rect 498198 0 498254 800
rect 499210 0 499266 800
rect 500222 0 500278 800
<< obsm2 >>
rect 480 601841 2078 601897
rect 2246 601841 6402 601897
rect 6570 601841 10818 601897
rect 10986 601841 15234 601897
rect 15402 601841 19650 601897
rect 19818 601841 23974 601897
rect 24142 601841 28390 601897
rect 28558 601841 32806 601897
rect 32974 601841 37222 601897
rect 37390 601841 41546 601897
rect 41714 601841 45962 601897
rect 46130 601841 50378 601897
rect 50546 601841 54794 601897
rect 54962 601841 59118 601897
rect 59286 601841 63534 601897
rect 63702 601841 67950 601897
rect 68118 601841 72366 601897
rect 72534 601841 76690 601897
rect 76858 601841 81106 601897
rect 81274 601841 85522 601897
rect 85690 601841 89938 601897
rect 90106 601841 94262 601897
rect 94430 601841 98678 601897
rect 98846 601841 103094 601897
rect 103262 601841 107510 601897
rect 107678 601841 111834 601897
rect 112002 601841 116250 601897
rect 116418 601841 120666 601897
rect 120834 601841 125082 601897
rect 125250 601841 129406 601897
rect 129574 601841 133822 601897
rect 133990 601841 138238 601897
rect 138406 601841 142654 601897
rect 142822 601841 146978 601897
rect 147146 601841 151394 601897
rect 151562 601841 155810 601897
rect 155978 601841 160226 601897
rect 160394 601841 164550 601897
rect 164718 601841 168966 601897
rect 169134 601841 173382 601897
rect 173550 601841 177798 601897
rect 177966 601841 182122 601897
rect 182290 601841 186538 601897
rect 186706 601841 190954 601897
rect 191122 601841 195370 601897
rect 195538 601841 199694 601897
rect 199862 601841 204110 601897
rect 204278 601841 208526 601897
rect 208694 601841 212942 601897
rect 213110 601841 217266 601897
rect 217434 601841 221682 601897
rect 221850 601841 226098 601897
rect 226266 601841 230514 601897
rect 230682 601841 234838 601897
rect 235006 601841 239254 601897
rect 239422 601841 243670 601897
rect 243838 601841 248086 601897
rect 248254 601841 252502 601897
rect 252670 601841 256826 601897
rect 256994 601841 261242 601897
rect 261410 601841 265658 601897
rect 265826 601841 270074 601897
rect 270242 601841 274398 601897
rect 274566 601841 278814 601897
rect 278982 601841 283230 601897
rect 283398 601841 287646 601897
rect 287814 601841 291970 601897
rect 292138 601841 296386 601897
rect 296554 601841 300802 601897
rect 300970 601841 305218 601897
rect 305386 601841 309542 601897
rect 309710 601841 313958 601897
rect 314126 601841 318374 601897
rect 318542 601841 322790 601897
rect 322958 601841 327114 601897
rect 327282 601841 331530 601897
rect 331698 601841 335946 601897
rect 336114 601841 340362 601897
rect 340530 601841 344686 601897
rect 344854 601841 349102 601897
rect 349270 601841 353518 601897
rect 353686 601841 357934 601897
rect 358102 601841 362258 601897
rect 362426 601841 366674 601897
rect 366842 601841 371090 601897
rect 371258 601841 375506 601897
rect 375674 601841 379830 601897
rect 379998 601841 384246 601897
rect 384414 601841 388662 601897
rect 388830 601841 393078 601897
rect 393246 601841 397402 601897
rect 397570 601841 401818 601897
rect 401986 601841 406234 601897
rect 406402 601841 410650 601897
rect 410818 601841 414974 601897
rect 415142 601841 419390 601897
rect 419558 601841 423806 601897
rect 423974 601841 428222 601897
rect 428390 601841 432546 601897
rect 432714 601841 436962 601897
rect 437130 601841 441378 601897
rect 441546 601841 445794 601897
rect 445962 601841 450118 601897
rect 450286 601841 454534 601897
rect 454702 601841 458950 601897
rect 459118 601841 463366 601897
rect 463534 601841 467690 601897
rect 467858 601841 472106 601897
rect 472274 601841 476522 601897
rect 476690 601841 480938 601897
rect 481106 601841 485262 601897
rect 485430 601841 489678 601897
rect 489846 601841 494094 601897
rect 494262 601841 498510 601897
rect 498678 601841 500276 601897
rect 480 856 500276 601841
rect 590 734 1434 856
rect 1602 734 2446 856
rect 2614 734 3458 856
rect 3626 734 4470 856
rect 4638 734 5482 856
rect 5650 734 6494 856
rect 6662 734 7506 856
rect 7674 734 8518 856
rect 8686 734 9530 856
rect 9698 734 10542 856
rect 10710 734 11554 856
rect 11722 734 12566 856
rect 12734 734 13578 856
rect 13746 734 14590 856
rect 14758 734 15602 856
rect 15770 734 16614 856
rect 16782 734 17626 856
rect 17794 734 18638 856
rect 18806 734 19650 856
rect 19818 734 20662 856
rect 20830 734 21674 856
rect 21842 734 22686 856
rect 22854 734 23698 856
rect 23866 734 24802 856
rect 24970 734 25814 856
rect 25982 734 26826 856
rect 26994 734 27838 856
rect 28006 734 28850 856
rect 29018 734 29862 856
rect 30030 734 30874 856
rect 31042 734 31886 856
rect 32054 734 32898 856
rect 33066 734 33910 856
rect 34078 734 34922 856
rect 35090 734 35934 856
rect 36102 734 36946 856
rect 37114 734 37958 856
rect 38126 734 38970 856
rect 39138 734 39982 856
rect 40150 734 40994 856
rect 41162 734 42006 856
rect 42174 734 43018 856
rect 43186 734 44030 856
rect 44198 734 45042 856
rect 45210 734 46054 856
rect 46222 734 47066 856
rect 47234 734 48170 856
rect 48338 734 49182 856
rect 49350 734 50194 856
rect 50362 734 51206 856
rect 51374 734 52218 856
rect 52386 734 53230 856
rect 53398 734 54242 856
rect 54410 734 55254 856
rect 55422 734 56266 856
rect 56434 734 57278 856
rect 57446 734 58290 856
rect 58458 734 59302 856
rect 59470 734 60314 856
rect 60482 734 61326 856
rect 61494 734 62338 856
rect 62506 734 63350 856
rect 63518 734 64362 856
rect 64530 734 65374 856
rect 65542 734 66386 856
rect 66554 734 67398 856
rect 67566 734 68410 856
rect 68578 734 69422 856
rect 69590 734 70434 856
rect 70602 734 71446 856
rect 71614 734 72550 856
rect 72718 734 73562 856
rect 73730 734 74574 856
rect 74742 734 75586 856
rect 75754 734 76598 856
rect 76766 734 77610 856
rect 77778 734 78622 856
rect 78790 734 79634 856
rect 79802 734 80646 856
rect 80814 734 81658 856
rect 81826 734 82670 856
rect 82838 734 83682 856
rect 83850 734 84694 856
rect 84862 734 85706 856
rect 85874 734 86718 856
rect 86886 734 87730 856
rect 87898 734 88742 856
rect 88910 734 89754 856
rect 89922 734 90766 856
rect 90934 734 91778 856
rect 91946 734 92790 856
rect 92958 734 93802 856
rect 93970 734 94814 856
rect 94982 734 95918 856
rect 96086 734 96930 856
rect 97098 734 97942 856
rect 98110 734 98954 856
rect 99122 734 99966 856
rect 100134 734 100978 856
rect 101146 734 101990 856
rect 102158 734 103002 856
rect 103170 734 104014 856
rect 104182 734 105026 856
rect 105194 734 106038 856
rect 106206 734 107050 856
rect 107218 734 108062 856
rect 108230 734 109074 856
rect 109242 734 110086 856
rect 110254 734 111098 856
rect 111266 734 112110 856
rect 112278 734 113122 856
rect 113290 734 114134 856
rect 114302 734 115146 856
rect 115314 734 116158 856
rect 116326 734 117170 856
rect 117338 734 118182 856
rect 118350 734 119194 856
rect 119362 734 120298 856
rect 120466 734 121310 856
rect 121478 734 122322 856
rect 122490 734 123334 856
rect 123502 734 124346 856
rect 124514 734 125358 856
rect 125526 734 126370 856
rect 126538 734 127382 856
rect 127550 734 128394 856
rect 128562 734 129406 856
rect 129574 734 130418 856
rect 130586 734 131430 856
rect 131598 734 132442 856
rect 132610 734 133454 856
rect 133622 734 134466 856
rect 134634 734 135478 856
rect 135646 734 136490 856
rect 136658 734 137502 856
rect 137670 734 138514 856
rect 138682 734 139526 856
rect 139694 734 140538 856
rect 140706 734 141550 856
rect 141718 734 142562 856
rect 142730 734 143666 856
rect 143834 734 144678 856
rect 144846 734 145690 856
rect 145858 734 146702 856
rect 146870 734 147714 856
rect 147882 734 148726 856
rect 148894 734 149738 856
rect 149906 734 150750 856
rect 150918 734 151762 856
rect 151930 734 152774 856
rect 152942 734 153786 856
rect 153954 734 154798 856
rect 154966 734 155810 856
rect 155978 734 156822 856
rect 156990 734 157834 856
rect 158002 734 158846 856
rect 159014 734 159858 856
rect 160026 734 160870 856
rect 161038 734 161882 856
rect 162050 734 162894 856
rect 163062 734 163906 856
rect 164074 734 164918 856
rect 165086 734 165930 856
rect 166098 734 166942 856
rect 167110 734 168046 856
rect 168214 734 169058 856
rect 169226 734 170070 856
rect 170238 734 171082 856
rect 171250 734 172094 856
rect 172262 734 173106 856
rect 173274 734 174118 856
rect 174286 734 175130 856
rect 175298 734 176142 856
rect 176310 734 177154 856
rect 177322 734 178166 856
rect 178334 734 179178 856
rect 179346 734 180190 856
rect 180358 734 181202 856
rect 181370 734 182214 856
rect 182382 734 183226 856
rect 183394 734 184238 856
rect 184406 734 185250 856
rect 185418 734 186262 856
rect 186430 734 187274 856
rect 187442 734 188286 856
rect 188454 734 189298 856
rect 189466 734 190310 856
rect 190478 734 191414 856
rect 191582 734 192426 856
rect 192594 734 193438 856
rect 193606 734 194450 856
rect 194618 734 195462 856
rect 195630 734 196474 856
rect 196642 734 197486 856
rect 197654 734 198498 856
rect 198666 734 199510 856
rect 199678 734 200522 856
rect 200690 734 201534 856
rect 201702 734 202546 856
rect 202714 734 203558 856
rect 203726 734 204570 856
rect 204738 734 205582 856
rect 205750 734 206594 856
rect 206762 734 207606 856
rect 207774 734 208618 856
rect 208786 734 209630 856
rect 209798 734 210642 856
rect 210810 734 211654 856
rect 211822 734 212666 856
rect 212834 734 213678 856
rect 213846 734 214690 856
rect 214858 734 215794 856
rect 215962 734 216806 856
rect 216974 734 217818 856
rect 217986 734 218830 856
rect 218998 734 219842 856
rect 220010 734 220854 856
rect 221022 734 221866 856
rect 222034 734 222878 856
rect 223046 734 223890 856
rect 224058 734 224902 856
rect 225070 734 225914 856
rect 226082 734 226926 856
rect 227094 734 227938 856
rect 228106 734 228950 856
rect 229118 734 229962 856
rect 230130 734 230974 856
rect 231142 734 231986 856
rect 232154 734 232998 856
rect 233166 734 234010 856
rect 234178 734 235022 856
rect 235190 734 236034 856
rect 236202 734 237046 856
rect 237214 734 238058 856
rect 238226 734 239162 856
rect 239330 734 240174 856
rect 240342 734 241186 856
rect 241354 734 242198 856
rect 242366 734 243210 856
rect 243378 734 244222 856
rect 244390 734 245234 856
rect 245402 734 246246 856
rect 246414 734 247258 856
rect 247426 734 248270 856
rect 248438 734 249282 856
rect 249450 734 250294 856
rect 250462 734 251306 856
rect 251474 734 252318 856
rect 252486 734 253330 856
rect 253498 734 254342 856
rect 254510 734 255354 856
rect 255522 734 256366 856
rect 256534 734 257378 856
rect 257546 734 258390 856
rect 258558 734 259402 856
rect 259570 734 260414 856
rect 260582 734 261426 856
rect 261594 734 262438 856
rect 262606 734 263542 856
rect 263710 734 264554 856
rect 264722 734 265566 856
rect 265734 734 266578 856
rect 266746 734 267590 856
rect 267758 734 268602 856
rect 268770 734 269614 856
rect 269782 734 270626 856
rect 270794 734 271638 856
rect 271806 734 272650 856
rect 272818 734 273662 856
rect 273830 734 274674 856
rect 274842 734 275686 856
rect 275854 734 276698 856
rect 276866 734 277710 856
rect 277878 734 278722 856
rect 278890 734 279734 856
rect 279902 734 280746 856
rect 280914 734 281758 856
rect 281926 734 282770 856
rect 282938 734 283782 856
rect 283950 734 284794 856
rect 284962 734 285806 856
rect 285974 734 286910 856
rect 287078 734 287922 856
rect 288090 734 288934 856
rect 289102 734 289946 856
rect 290114 734 290958 856
rect 291126 734 291970 856
rect 292138 734 292982 856
rect 293150 734 293994 856
rect 294162 734 295006 856
rect 295174 734 296018 856
rect 296186 734 297030 856
rect 297198 734 298042 856
rect 298210 734 299054 856
rect 299222 734 300066 856
rect 300234 734 301078 856
rect 301246 734 302090 856
rect 302258 734 303102 856
rect 303270 734 304114 856
rect 304282 734 305126 856
rect 305294 734 306138 856
rect 306306 734 307150 856
rect 307318 734 308162 856
rect 308330 734 309174 856
rect 309342 734 310186 856
rect 310354 734 311290 856
rect 311458 734 312302 856
rect 312470 734 313314 856
rect 313482 734 314326 856
rect 314494 734 315338 856
rect 315506 734 316350 856
rect 316518 734 317362 856
rect 317530 734 318374 856
rect 318542 734 319386 856
rect 319554 734 320398 856
rect 320566 734 321410 856
rect 321578 734 322422 856
rect 322590 734 323434 856
rect 323602 734 324446 856
rect 324614 734 325458 856
rect 325626 734 326470 856
rect 326638 734 327482 856
rect 327650 734 328494 856
rect 328662 734 329506 856
rect 329674 734 330518 856
rect 330686 734 331530 856
rect 331698 734 332542 856
rect 332710 734 333554 856
rect 333722 734 334658 856
rect 334826 734 335670 856
rect 335838 734 336682 856
rect 336850 734 337694 856
rect 337862 734 338706 856
rect 338874 734 339718 856
rect 339886 734 340730 856
rect 340898 734 341742 856
rect 341910 734 342754 856
rect 342922 734 343766 856
rect 343934 734 344778 856
rect 344946 734 345790 856
rect 345958 734 346802 856
rect 346970 734 347814 856
rect 347982 734 348826 856
rect 348994 734 349838 856
rect 350006 734 350850 856
rect 351018 734 351862 856
rect 352030 734 352874 856
rect 353042 734 353886 856
rect 354054 734 354898 856
rect 355066 734 355910 856
rect 356078 734 356922 856
rect 357090 734 357934 856
rect 358102 734 359038 856
rect 359206 734 360050 856
rect 360218 734 361062 856
rect 361230 734 362074 856
rect 362242 734 363086 856
rect 363254 734 364098 856
rect 364266 734 365110 856
rect 365278 734 366122 856
rect 366290 734 367134 856
rect 367302 734 368146 856
rect 368314 734 369158 856
rect 369326 734 370170 856
rect 370338 734 371182 856
rect 371350 734 372194 856
rect 372362 734 373206 856
rect 373374 734 374218 856
rect 374386 734 375230 856
rect 375398 734 376242 856
rect 376410 734 377254 856
rect 377422 734 378266 856
rect 378434 734 379278 856
rect 379446 734 380290 856
rect 380458 734 381302 856
rect 381470 734 382406 856
rect 382574 734 383418 856
rect 383586 734 384430 856
rect 384598 734 385442 856
rect 385610 734 386454 856
rect 386622 734 387466 856
rect 387634 734 388478 856
rect 388646 734 389490 856
rect 389658 734 390502 856
rect 390670 734 391514 856
rect 391682 734 392526 856
rect 392694 734 393538 856
rect 393706 734 394550 856
rect 394718 734 395562 856
rect 395730 734 396574 856
rect 396742 734 397586 856
rect 397754 734 398598 856
rect 398766 734 399610 856
rect 399778 734 400622 856
rect 400790 734 401634 856
rect 401802 734 402646 856
rect 402814 734 403658 856
rect 403826 734 404670 856
rect 404838 734 405682 856
rect 405850 734 406786 856
rect 406954 734 407798 856
rect 407966 734 408810 856
rect 408978 734 409822 856
rect 409990 734 410834 856
rect 411002 734 411846 856
rect 412014 734 412858 856
rect 413026 734 413870 856
rect 414038 734 414882 856
rect 415050 734 415894 856
rect 416062 734 416906 856
rect 417074 734 417918 856
rect 418086 734 418930 856
rect 419098 734 419942 856
rect 420110 734 420954 856
rect 421122 734 421966 856
rect 422134 734 422978 856
rect 423146 734 423990 856
rect 424158 734 425002 856
rect 425170 734 426014 856
rect 426182 734 427026 856
rect 427194 734 428038 856
rect 428206 734 429050 856
rect 429218 734 430154 856
rect 430322 734 431166 856
rect 431334 734 432178 856
rect 432346 734 433190 856
rect 433358 734 434202 856
rect 434370 734 435214 856
rect 435382 734 436226 856
rect 436394 734 437238 856
rect 437406 734 438250 856
rect 438418 734 439262 856
rect 439430 734 440274 856
rect 440442 734 441286 856
rect 441454 734 442298 856
rect 442466 734 443310 856
rect 443478 734 444322 856
rect 444490 734 445334 856
rect 445502 734 446346 856
rect 446514 734 447358 856
rect 447526 734 448370 856
rect 448538 734 449382 856
rect 449550 734 450394 856
rect 450562 734 451406 856
rect 451574 734 452418 856
rect 452586 734 453430 856
rect 453598 734 454534 856
rect 454702 734 455546 856
rect 455714 734 456558 856
rect 456726 734 457570 856
rect 457738 734 458582 856
rect 458750 734 459594 856
rect 459762 734 460606 856
rect 460774 734 461618 856
rect 461786 734 462630 856
rect 462798 734 463642 856
rect 463810 734 464654 856
rect 464822 734 465666 856
rect 465834 734 466678 856
rect 466846 734 467690 856
rect 467858 734 468702 856
rect 468870 734 469714 856
rect 469882 734 470726 856
rect 470894 734 471738 856
rect 471906 734 472750 856
rect 472918 734 473762 856
rect 473930 734 474774 856
rect 474942 734 475786 856
rect 475954 734 476798 856
rect 476966 734 477902 856
rect 478070 734 478914 856
rect 479082 734 479926 856
rect 480094 734 480938 856
rect 481106 734 481950 856
rect 482118 734 482962 856
rect 483130 734 483974 856
rect 484142 734 484986 856
rect 485154 734 485998 856
rect 486166 734 487010 856
rect 487178 734 488022 856
rect 488190 734 489034 856
rect 489202 734 490046 856
rect 490214 734 491058 856
rect 491226 734 492070 856
rect 492238 734 493082 856
rect 493250 734 494094 856
rect 494262 734 495106 856
rect 495274 734 496118 856
rect 496286 734 497130 856
rect 497298 734 498142 856
rect 498310 734 499154 856
rect 499322 734 500166 856
<< obsm3 >>
rect 3233 2143 496048 600065
<< metal4 >>
rect 4208 2128 4528 600080
rect 19568 2128 19888 600080
rect 34928 2128 35248 600080
rect 50288 2128 50608 600080
rect 65648 2128 65968 600080
rect 81008 2128 81328 600080
rect 96368 2128 96688 600080
rect 111728 2128 112048 600080
rect 127088 2128 127408 600080
rect 142448 2128 142768 600080
rect 157808 2128 158128 600080
rect 173168 2128 173488 600080
rect 188528 2128 188848 600080
rect 203888 2128 204208 600080
rect 219248 2128 219568 600080
rect 234608 2128 234928 600080
rect 249968 2128 250288 600080
rect 265328 2128 265648 600080
rect 280688 2128 281008 600080
rect 296048 2128 296368 600080
rect 311408 2128 311728 600080
rect 326768 2128 327088 600080
rect 342128 2128 342448 600080
rect 357488 2128 357808 600080
rect 372848 2128 373168 600080
rect 388208 2128 388528 600080
rect 403568 2128 403888 600080
rect 418928 2128 419248 600080
rect 434288 2128 434608 600080
rect 449648 2128 449968 600080
rect 465008 2128 465328 600080
rect 480368 2128 480688 600080
rect 495728 2128 496048 600080
<< obsm4 >>
rect 19379 109787 19488 538797
rect 19968 109787 34848 538797
rect 35328 109787 50208 538797
rect 50688 109787 65568 538797
rect 66048 109787 80928 538797
rect 81408 109787 96288 538797
rect 96768 109787 111648 538797
rect 112128 109787 127008 538797
rect 127488 109787 142368 538797
rect 142848 109787 157728 538797
rect 158208 109787 173088 538797
rect 173568 109787 188448 538797
rect 188928 109787 203808 538797
rect 204288 109787 219168 538797
rect 219648 109787 234528 538797
rect 235008 109787 249888 538797
rect 250368 109787 265248 538797
rect 265728 109787 280608 538797
rect 281088 109787 295968 538797
rect 296448 109787 311328 538797
rect 311808 109787 326688 538797
rect 327168 109787 342048 538797
rect 342528 109787 357408 538797
rect 357888 109787 372768 538797
rect 373248 109787 388128 538797
rect 388608 109787 403488 538797
rect 403968 109787 418848 538797
rect 419328 109787 434208 538797
rect 434688 109787 448533 538797
<< labels >>
rlabel metal2 s 2134 601897 2190 602697 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 133878 601897 133934 602697 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 147034 601897 147090 602697 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 160282 601897 160338 602697 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 173438 601897 173494 602697 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 186594 601897 186650 602697 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 199750 601897 199806 602697 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 212998 601897 213054 602697 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 226154 601897 226210 602697 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 239310 601897 239366 602697 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 252558 601897 252614 602697 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 15290 601897 15346 602697 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 265714 601897 265770 602697 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 278870 601897 278926 602697 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 292026 601897 292082 602697 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 305274 601897 305330 602697 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 318430 601897 318486 602697 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 331586 601897 331642 602697 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 344742 601897 344798 602697 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 357990 601897 358046 602697 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 371146 601897 371202 602697 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 384302 601897 384358 602697 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 28446 601897 28502 602697 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 397458 601897 397514 602697 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 410706 601897 410762 602697 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 423862 601897 423918 602697 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 437018 601897 437074 602697 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 450174 601897 450230 602697 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 463422 601897 463478 602697 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 476578 601897 476634 602697 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 489734 601897 489790 602697 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 41602 601897 41658 602697 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 54850 601897 54906 602697 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 68006 601897 68062 602697 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 81162 601897 81218 602697 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 94318 601897 94374 602697 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 107566 601897 107622 602697 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 120722 601897 120778 602697 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6458 601897 6514 602697 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 138294 601897 138350 602697 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 151450 601897 151506 602697 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 164606 601897 164662 602697 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 177854 601897 177910 602697 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 191010 601897 191066 602697 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 204166 601897 204222 602697 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 217322 601897 217378 602697 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 230570 601897 230626 602697 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 243726 601897 243782 602697 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 256882 601897 256938 602697 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 19706 601897 19762 602697 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 270130 601897 270186 602697 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 283286 601897 283342 602697 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 296442 601897 296498 602697 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 309598 601897 309654 602697 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 322846 601897 322902 602697 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 336002 601897 336058 602697 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 349158 601897 349214 602697 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 362314 601897 362370 602697 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 375562 601897 375618 602697 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 388718 601897 388774 602697 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 32862 601897 32918 602697 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 401874 601897 401930 602697 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 415030 601897 415086 602697 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 428278 601897 428334 602697 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 441434 601897 441490 602697 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 454590 601897 454646 602697 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 467746 601897 467802 602697 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 480994 601897 481050 602697 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 494150 601897 494206 602697 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 46018 601897 46074 602697 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 59174 601897 59230 602697 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 72422 601897 72478 602697 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 85578 601897 85634 602697 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 98734 601897 98790 602697 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 111890 601897 111946 602697 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 125138 601897 125194 602697 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 10874 601897 10930 602697 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 142710 601897 142766 602697 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 155866 601897 155922 602697 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 169022 601897 169078 602697 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 182178 601897 182234 602697 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 195426 601897 195482 602697 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 208582 601897 208638 602697 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 221738 601897 221794 602697 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 234894 601897 234950 602697 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 248142 601897 248198 602697 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 261298 601897 261354 602697 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 24030 601897 24086 602697 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 274454 601897 274510 602697 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 287702 601897 287758 602697 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 300858 601897 300914 602697 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 314014 601897 314070 602697 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 327170 601897 327226 602697 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 340418 601897 340474 602697 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 353574 601897 353630 602697 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 366730 601897 366786 602697 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 379886 601897 379942 602697 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 393134 601897 393190 602697 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 37278 601897 37334 602697 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 406290 601897 406346 602697 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 419446 601897 419502 602697 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 432602 601897 432658 602697 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 445850 601897 445906 602697 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 459006 601897 459062 602697 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 472162 601897 472218 602697 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 485318 601897 485374 602697 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 498566 601897 498622 602697 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 50434 601897 50490 602697 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 63590 601897 63646 602697 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 76746 601897 76802 602697 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 89994 601897 90050 602697 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 103150 601897 103206 602697 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 116306 601897 116362 602697 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 129462 601897 129518 602697 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 498198 0 498254 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 499210 0 499266 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 500222 0 500278 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 412914 0 412970 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 415950 0 416006 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 418986 0 419042 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 422022 0 422078 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 425058 0 425114 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 428094 0 428150 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 431222 0 431278 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 434258 0 434314 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 437294 0 437350 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 440330 0 440386 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 443366 0 443422 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 446402 0 446458 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 449438 0 449494 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 452474 0 452530 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 455602 0 455658 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 458638 0 458694 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 461674 0 461730 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 464710 0 464766 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 467746 0 467802 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 470782 0 470838 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 473818 0 473874 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 476854 0 476910 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 479982 0 480038 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 483018 0 483074 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 486054 0 486110 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 489090 0 489146 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 492126 0 492182 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 495162 0 495218 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 181258 0 181314 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 184294 0 184350 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 187330 0 187386 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 190366 0 190422 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 199566 0 199622 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 214746 0 214802 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 217874 0 217930 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 220910 0 220966 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 223946 0 224002 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 226982 0 227038 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 233054 0 233110 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 236090 0 236146 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 239218 0 239274 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 242254 0 242310 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 245290 0 245346 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 248326 0 248382 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 251362 0 251418 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 257434 0 257490 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 260470 0 260526 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 272706 0 272762 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 278778 0 278834 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 281814 0 281870 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 284850 0 284906 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 287978 0 288034 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 291014 0 291070 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 294050 0 294106 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 297086 0 297142 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 300122 0 300178 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 303158 0 303214 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 306194 0 306250 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 309230 0 309286 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 312358 0 312414 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 315394 0 315450 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 318430 0 318486 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 321466 0 321522 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 324502 0 324558 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 327538 0 327594 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 330574 0 330630 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 333610 0 333666 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 336738 0 336794 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 339774 0 339830 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 342810 0 342866 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 345846 0 345902 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 348882 0 348938 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 351918 0 351974 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 354954 0 355010 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 357990 0 358046 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 361118 0 361174 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 364154 0 364210 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 367190 0 367246 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 370226 0 370282 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 373262 0 373318 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 376298 0 376354 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 379334 0 379390 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 382462 0 382518 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 385498 0 385554 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 388534 0 388590 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 391570 0 391626 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 394606 0 394662 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 397642 0 397698 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 400678 0 400734 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 403714 0 403770 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 406842 0 406898 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 409878 0 409934 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 413926 0 413982 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 416962 0 417018 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 419998 0 420054 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 423034 0 423090 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 426070 0 426126 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 429106 0 429162 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 432234 0 432290 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 435270 0 435326 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 438306 0 438362 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 441342 0 441398 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 444378 0 444434 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 447414 0 447470 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 450450 0 450506 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 453486 0 453542 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 456614 0 456670 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 459650 0 459706 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 462686 0 462742 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 465722 0 465778 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 468758 0 468814 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 471794 0 471850 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 474830 0 474886 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 477958 0 478014 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 480994 0 481050 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 484030 0 484086 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 487066 0 487122 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 490102 0 490158 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 493138 0 493194 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 496174 0 496230 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 154854 0 154910 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 157890 0 157946 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 160926 0 160982 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 166998 0 167054 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 170126 0 170182 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 176198 0 176254 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 179234 0 179290 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 182270 0 182326 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 185306 0 185362 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 188342 0 188398 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 191470 0 191526 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 194506 0 194562 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 197542 0 197598 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 200578 0 200634 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 203614 0 203670 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 206650 0 206706 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 209686 0 209742 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 212722 0 212778 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 215850 0 215906 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 218886 0 218942 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 221922 0 221978 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 224958 0 225014 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 227994 0 228050 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 231030 0 231086 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 234066 0 234122 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 237102 0 237158 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 240230 0 240286 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 243266 0 243322 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 246302 0 246358 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 249338 0 249394 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 252374 0 252430 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 255410 0 255466 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 258446 0 258502 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 261482 0 261538 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 264610 0 264666 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 267646 0 267702 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 270682 0 270738 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 273718 0 273774 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 276754 0 276810 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 279790 0 279846 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 282826 0 282882 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 285862 0 285918 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 288990 0 289046 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 292026 0 292082 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 295062 0 295118 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 298098 0 298154 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 301134 0 301190 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 304170 0 304226 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 307206 0 307262 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 310242 0 310298 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 313370 0 313426 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 316406 0 316462 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 319442 0 319498 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 322478 0 322534 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 325514 0 325570 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 328550 0 328606 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 331586 0 331642 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 334714 0 334770 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 337750 0 337806 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 340786 0 340842 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 343822 0 343878 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 346858 0 346914 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 349894 0 349950 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 352930 0 352986 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 355966 0 356022 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 359094 0 359150 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 362130 0 362186 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 365166 0 365222 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 368202 0 368258 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 371238 0 371294 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 374274 0 374330 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 377310 0 377366 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 380346 0 380402 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 133510 0 133566 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 383474 0 383530 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 386510 0 386566 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 389546 0 389602 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 392582 0 392638 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 395618 0 395674 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 398654 0 398710 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 401690 0 401746 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 404726 0 404782 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 407854 0 407910 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 410890 0 410946 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 414938 0 414994 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 417974 0 418030 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 421010 0 421066 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 424046 0 424102 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 427082 0 427138 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 430210 0 430266 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 433246 0 433302 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 436282 0 436338 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 439318 0 439374 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 442354 0 442410 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 445390 0 445446 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 448426 0 448482 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 451462 0 451518 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 454590 0 454646 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 457626 0 457682 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 460662 0 460718 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 463698 0 463754 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 466734 0 466790 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 469770 0 469826 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 472806 0 472862 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 475842 0 475898 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 478970 0 479026 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 482006 0 482062 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 485042 0 485098 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 488078 0 488134 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 491114 0 491170 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 494150 0 494206 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 497186 0 497242 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 180246 0 180302 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 201590 0 201646 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 210698 0 210754 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 213734 0 213790 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 216862 0 216918 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 222934 0 222990 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 229006 0 229062 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 232042 0 232098 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 238114 0 238170 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 244278 0 244334 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 250350 0 250406 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 256422 0 256478 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 259458 0 259514 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 262494 0 262550 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 265622 0 265678 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 268658 0 268714 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 271694 0 271750 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 274730 0 274786 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 277766 0 277822 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 280802 0 280858 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 283838 0 283894 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 286966 0 287022 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 290002 0 290058 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 293038 0 293094 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 296074 0 296130 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 299110 0 299166 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 302146 0 302202 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 305182 0 305238 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 308218 0 308274 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 311346 0 311402 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 314382 0 314438 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 317418 0 317474 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 320454 0 320510 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 323490 0 323546 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 326526 0 326582 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 329562 0 329618 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 332598 0 332654 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 335726 0 335782 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 338762 0 338818 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 341798 0 341854 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 344834 0 344890 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 347870 0 347926 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 350906 0 350962 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 353942 0 353998 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 356978 0 357034 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 360106 0 360162 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 363142 0 363198 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 366178 0 366234 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 369214 0 369270 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 372250 0 372306 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 375286 0 375342 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 378322 0 378378 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 381358 0 381414 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 384486 0 384542 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 387522 0 387578 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 390558 0 390614 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 393594 0 393650 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 396630 0 396686 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 399666 0 399722 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 402702 0 402758 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 405738 0 405794 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 408866 0 408922 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 411902 0 411958 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 434288 2128 434608 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 465008 2128 465328 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 495728 2128 496048 600080 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 418928 2128 419248 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 449648 2128 449968 600080 6 vssd1
port 503 nsew ground input
rlabel metal4 s 480368 2128 480688 600080 6 vssd1
port 503 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 500829 602697
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 361836910
string GDS_START 1169594
<< end >>

